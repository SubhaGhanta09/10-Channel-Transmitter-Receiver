PK   �|�X_�ά9=  m8    cirkitFile.json�o�6������.:���ٹ�@23��̤�dg.�%Q�sǱ{��yl�t���M�����q�JgwӘ�m�*},��,�,�|z��W��M��>��n��N_�9;}n��ӣ������b{}��Mx�������j�ӛX571t�u��"6������+]����UյF�t|w!.��˯�9{�@K�f�J2Ix�������U��^4��m]U7^TZ�X�Z�ʶ�p����p�Oq���[��ŅBk_a�_��D��S<��i@�
�[{ � V�^"k_#k�=���B�koc�mL����٪鄮��Ѻ���(t�����F ��och'�j�K�{�VΛPE�H�j��ѵ�h���M�5����t�n�ʫZVA[����h|�w����
��謪B/�J��UA馲��ާ6���� ��*������:����Gr^W��Qic��_�����A�'b�WB���BHO@�܁�[��w��{|���7�?ě�&l.�\���7��O��[�7 �`&�h��`�j�z�����kd�zŊH5�+"Q8<VD��w_h)��wBh�ߓ�E$
|w��(�!ZD���a��D�u|��(�-"Q�}'ZD���N��D���h�B�}'ZD���N��D���h���m�w*��D�Hx߉�(�-"Q�}'ZD���N��D���h�B�}'ZD���N��D���h��;�"�����O
�k���xϋ�(�-"Q�=/Z��gU��T��o�E$
��F�Hx��1|��Y�6� �u�{}��D�1�E$
��F���#?+c�
����E$
�x-"=�x���(�~-"Q���D��ODb����WD�� 6���͟A����T}�7����_�)I�V� (��Lܮb8=%ݞ8<��-��������#�Z:q�hu�huGJ�t)�՝��)�ҥ�KIU4U
�C�����CMtB&���lI���ö�-i�"l�MtB&����+�K�m���ŊH�-6�	�8�s%-V4��b��ŊH�-6�	�8��%-V4��b��ŊH�-6�	�8�H�(8.�b�m2(���P�m6�
�<�V���#d��8F� ��dZ> �Nfǽ���ā��zt�H�Okq�M��|�kH�w j~֒���C�i���"�员/q K˗�v�4nb> �˫R��GE1���4��#�i�����J �O4���1_^�D�?�臖���꫒��(� 6旓���(ؘ�:y$�F�qRM�|@̗���8h��b��B�X�Q�1_^�H�?⨇����Lb�G=�|@̗ד�8��b���X�Q-��5�ē���Z> �˫���G���1_^7M�?�o>�|@̗W|�zv$��H��C��8���b��ʞX��-��� ��#�?h���/g6 �q�A��|9'����Z> ���$��G��1_΃A�?M��1_��A�?������r�b���|@̗���8���b���X�+���h��8����-��,9��#�?h���/��!�q�A��|93����Z> ��9���G��1_��D�?C��1_�DE�?������r-b���|@̗��8���b��y�X��-��i��#�?h���/g{#�q�A��|9O����Z> ��9��G��1_��G�?������r^BZ�Y������rFEb���|@̗sA�8���#|O��H����d�j�E窦�P���������=���q&ϕ��Sp��|��x���t�+/�	^y�8����ǹuW^>N����q6۵f�5;��Mv�\{=��&���i{�} �^�����{k�G��d����c���&�í�i���^����.hk�G��d籵��&�}����"�o�7����pI/no��\
����]��;&��v�Xys�����\�n.F�@��9n���9��-�樚/{q����WZu]�$&/ Z��n�́إ��e�}�ҡ`�R2]��J�ZD���݋.?t�F��䔺}Wi״U�I��oT���p���/�=�Vh��"�J�K+��j!C�A��._��SF�N�Uy�S�I�T �+[g}s��E�/߽�N(��ֆX��S/�4VW������&�{���=#c�U# )��d6���Z�gP{c�C�^r����6�>��b+ ]n�*�VV.�e�5�;T��˗�^���U��}u2t2��>���g���f�Ʃ�.i����d$�RD�m�z�慉�qj�%R�|��d�A�H��n^�/��q~_
�EƩ�(�&��Qga�t�"\I�f�'#Yn�"t����fB�����Havx2��)"A�,�݊����Z��(�IS�F��9�M��#�EVn!���0w^��;��ھ�U�GF�l��
�o�¦D�Ya�/í/��������˟1/x�m������aK"A"����,	�QqD����m ���� ��G�����M^��4Pn}�#2;"�+�#�;A��-�h'��5��΂LRw�#5�s�Vs;��w8�A��Zۀ#�T�=���!ɜ��$�@2ѹ�AR�M��z�dL�$�M�P��sG����LD��&m��{��u��?�H&C�d��D$IV���$�a�$1L�!b"�$��:4LT��0���n�M�ǩ$�a���d~�J�&T1��qI�ǩ$�a���d~�J�&�1��qE�ǩ$�a"�Wd~�J�&�1��qE�ǩ$�ab"�Wd~�JR�QI�D������s)�1��qM�ǩ$�dLd~\��q*I97��t/����6T/X5��d~�JR��E�D��5����sRQ}B�d~ܐ�q*I9w�7d~�JR��C��̐�qC�ǩ$�\4dLd~ܐ�q*I9g
�g`2?n��8���ۃ��̏[2?N%)� c"��̏/IB�Ԛ�扞�6��p}މ)+^0�J��q�r�d���
,��b�ʄ\*�^9X��U\�S,�K%�++�����E���4�`��6�~k����ߚ�R�u�J��q�F��6��u�J��)+�^�)i�:N�H��)+�^��z�v���8�#�^��z��R�u��F��ď4z��R�u�J2��	���4�4;CK0�\LAS��v��]�xO��B<�y�9�O���fh��R�' ���xh����Da,�0GK���f_,���b,�y-�n9"�ڼ��G�Q��m^ã[�Hxh��6������� -���J<���Xh��v�}�(v�%��В�'.�<�$O\�B<�y�ny�2Z��k�xt�� -���5�<���Xh��6����-O\�B<�y�(�ny�2Z��k]yt����m^��31�'.c�ڼ��G�<q-���5�<���^�B<�y-8�n�f+2MW��O\�x�2Z��k�yt����m�1��[����xhs����e,��C�s>��'.c�ڜ��G�<q-���,��<q-���\"<���Xh��6�D��-O\�B<�9��ny�2Z��9jxt˴��i)O\�y�2����m�ģ[����xhs�#���e,��C�s8��'.c�ڜ��G�<q-���Z,�5<q-����`<���Xh��6�8��-O\�B<�9W�ny�2Z��9�xt����mΝǣ[����xhs@���e,��C�s��'.c�ڜ��G�<q-���ܒ<���Xh��6��dѭ��Xh��6����-O\�B<�9g)�ny�2Z(�}��4M��J�>I���VC�:ƶ3Іni�RrӮ���Mv���<�+�,d�^)e!W�J)٭WJY�G�R�B�Rr>��:"㥱ޥ�c׊��ߥ�U׊���L׊���mB׊����8׊!��4V��K�Z14V���Z14V����Z14V�����^�Ɗ�v\+�h(Ac�K��sԊ�Њ޶��/*�U�\�ue�^8_��E؍��YVJ�i��a��]3��FH�k%�+��24��B���r�_V4B"��M�m ���~F4�F%D���V]W%���D�u�{�9!I9�\{�C�t(�T#�d��J�ZD����HJK#zo�j��*횶
2e�oT���P�R �(K���b%ET�N*��%�BU�I9�┑�uC�&7SKK�T �+[g}s��H�Q�6:�LRlb��$癔ZW��.�mo{��I9n/������RK�du���Z��^{c�{)�r��oC��*���T���r1�(��i\�^��e1��ִ�+R��۾�N��6)9�������H����H�����%)��1�6&R���٪鄮��Ѻ��ڨ�5*�r�FER���r�O@h'���^�k+�M��o��V����kT$�h���5RQk楨Ts��(�Uz�BHRڤ&[�J��\���I9Z�")C���ݩv^���YU�^&�W���&������kT$�h���܍��4Z������:�8���/^W��Qic���x����Q���F�6�^�b�pMv��Z�SO⤩\#m2`o��(����Q�L+Z�H�P#)ȅ�nz\R-bSI�=l��bo��N��F�m,x���n�IR#�D��b.���۰��/~�~˴����v{.���1�H��NBD$HmHBD$H�@BD$H1&	� 1ī$DD����	CMBD$H_aH����	� ��:D�"�6��&��@温$��G0&2�dΛJ��}��a"��@���$�݇C&2dN�J��}Ҥa"��̏SI���4Lt�o�8��d~�J��}S�a"��̏SI���4Ld~\��q*Ib����̏K2?N%I�fЄ�d~\��q*Ib7w����M
ݫ2?���8�$���A�D������s�1��qE�ǩ$�odLd~\��q*I9���d~�JR�aE�D�N��8��d~�JR�5D�D��5����sې1��qM�ǩ$�\*d�~���!��T�r�2&2?n��8���+�����&��M2?n��8�������̏2?N%)�!'c"��̏SI�k�ɘ���%��K�֯?��o���[&L XX��U\LֶSK%�++����ɺvj��z�`Vq1�5F-�P����.�NҌ�h��XX�8�E��c$�`�4Fa��$��8X��U\Lr�QK%�++����I^1j��z�`Vq1�)F-�P�����<-����<�e����.��x/���Xh��6�5��-O��B<�y�<�ny"0Z��s�yt����m^���[�H��xh�Z��Dc,��C�ה��'"c�ڼ6�G�<Q-���5><x�2Z��k�xt����m^sţ[�/bL��x�2��I����xh�8���e,��C�����'.c�ڼ&�G�<q-��浕<���Xh��6���-O\�B<�y�+�ny�2Z��kvy&&��e,��C����'.c�ڼ��G�<q-����<�e���4]�'.S<q���Xh��6����-O\�B<�9� �ny�2Z�͹xt����m����[����xhs�
���e,��C�sp��V��e,��C�s���'.c�ڜ�G�<q-����.<���Xh��6���-�J2��d<q���4O\�B<�9g�ny�2Z�͹�xt����m��ģ[����xhs.*���e,��C�sj�����e,��C�s���'.c�ڜ�G�<q-���\m<���Xh��6���-O\�B<�9w�n��|0�����O\fx�2Z�͹yt����m��ȣ[����xhsnI���e,��C�sd�����e,��C�s}��'.c�ڜ��G�<q-��>ݠ\��W]%��Zt�jZU����@��}�WJY�M�R�B6ٕR�x����y{���\�+�,d�^)e!�J)�WJY����ꈌ��z�6}]+��~��V]+�Ƃ�60]+�Ɔ��	]+�Ɗ�6�\+���X��.�k��X��^�k��X�Ҏ�k��X�Ҿ�k{]+^�=p����/m��V�Q+nB+zۺ�n���V�r�֕m{�|[����H��v*�r����m�")G�H
Mu4ER������WZu]�'���Q�]渽I9j/��Ї.
6�H)���R�B'�/`)�R�҈��Z�J����LAx�dtu�sT$�(K���b%ET�N*��!C�ADqER��8e��D]�P��M����5�3���Y�g)�r���N(�ۆX')�y&�֕�}��ބ�,ER��K4F� �F@ҩ���d-*��L�����R"�(K߆��Ul$)���me�bQ6]Ӹ�I9�bz�iuV�nM�}�U���mRrM���,ERhX��G��1�6&R���٪鄮��Ѻ��ڨ�5*�r�FER�֨��m��^�Kz񮭜7�����[�JW`�ER
��)Gk�R�!���V�9
!Ii��l�*��s]��kT$�h���V��UU�e�qUP��l��O����g�HJ���@����0���N'N���U�dT�+dAo_$�x�V"�h����M��j�N=���r��ɀ�MO�#��I9�52�"6����6��.����t�id�Ƃ'�H
�Q�Iy�r�~�1����뛋M���K��N���ۋ7�����������7�/��
��@�s�s��P�Y�0(�e���;ށB6�:��g�$�����; �n�17OV�����ws���B�\�nn��o�BG��]�Pu>E�ڥ�]+C��C��ڶ6�a1��_��ݽ���'�Y���û�l�1}>�	Y+�z:�M��z}� (�8lˍ�q �c �%�~T`�.�.˽�sj����w�!�ɯx��:�.�5��·(_DR��E�H
�8�H�"��&��	yE$��Q$e1V�CO����_�Q=<H
_4R=<H
_�S=<H
_�S=<H
?�P=<H
�-T�
��^�k_������踻� ��Q�����7��n�wFG���k+�VN������tc����k����;���|���Y!�h�_AP��l\[�%��dp���츉�]��p��}��*1�¿�����?������������7�����9������o�#:��t|��?���_����x�wv<�s�����_����z����|�3>�,��`V�O�M-����s\���H��@0O��)�Nk��O�3�?h���?��+�=�PP=�D
A�Z��/��_$���<���f�Bj�ݪi�@nU�[���mܮ�z;�
�טH^����u'.�f
��|� ���x'30�������|̃@�bZ&�󌟝y�]L��?f�s5��M�cF<s��O��?f��8��tN�cF0��dL��?Ms<�����h�3>�?�� ï1�sy�[(a���s/8��|T< rZ*�xv*�z�j":M�������6l��ˇ���~w������Mw��g̫�����|�E�!_
�-B�V��?�L���W�
�)5�¾W�C�E�!��^;�d"���N$��H�Ϛ���#��D��l覌��X�DY�ҹ#�
?�B 8�A��A���)����X�N ��f\86bBw,b�]�-�� f�6r�� �e	ԃ�!v�`9�2�n�,Z���X��@��-�xb�g��b8N�|�2�n�,�{��/C����r�SI�O�2�n�
,�?��/C����r�SE�O�2�n�,�?U�/C���r�SE�O�2�n,�?U�/#q�S���A�O�2�?��y&�5�?��/#q�S���A�O�2�k`���?��&p�����e$����8�+^�0)��}�&����e$o���8�-^ư����!p�����e�����x[��a	�WI�k�/^F� ��eKX�xy[{ok	��Tzj��3�&��:~$����(m��] �ۓG��|@�'.$��$��h���O\(b�)b���1_
]�����G��|���i����]��1�Gjw��Ԯ=�]d�4{D�5Nz�v'�H��G�+���j��1�Gjw��Ԯ;�]��^��E��)=R�\�v��Ү��h��aJ���;
?4���?�_d�4�����&���<r"��c'���:z"&j�i��Ó�q�iTJQ�9��fIT5�~�`���ǡ���XІ#�i̒:`"&��ީuHu 5!P�9��:��-���	�zj�F@MԄy���w��	��0���!uCLԄ�m.&#�M+&�Q/�`��a�GR$��A1!P�C�:�j�	��0�z��!m� Ԅ@M�WlQ�:�!&j¼ڌZ��Q1!P�r�:��b�	��0���!uCLԄy�"��(���	��JjRG1Ą@M�W�R��[1!P�U��:$��F>��:NQ�q���S�	��0�&��!u�BLԄy%4���bB�&̫��uH�5a^�N�C�8���	��yjR�)Ą@M�W��PS�)Ą@M��P�:N!&jq�Z��q
1!P�l�:��S�	��0g���!���7�q���S4u�BLԄ9����bB�&��P�uH�5aN�B�C�8���	sjR�)Ą@M�s���P�)Ą@M���P�:N!&j��Z��q
1!P�<K�:��S�	��0'���!u�BLԄ9����bB�&�ɸ�uH�5aN$F�C�8���	s�3jR�)Ą@M�3�Q�:N!&jm�X��:N!&j)�Z��q
1!P�,�:��S�	���m��iz�U2�ڬE窦�P��������n}���I�ƕ�O2,��~�xv�����+��$z]y�$A���'�TW^?ɀ���I�ҵ��6@�Nw�[+ k����
�Z�tS���v8�m� �%N7[+ ���8ݣk� �%Nw�Z+ k��}��
�Z�t秵}��{-���8ݖh���؄V��uU�xQi�b�j�+����:�.�6?�Ty���֮�+�W��ٗ[#ĩ�8����B��n�5B�̆�!����Q	Qy�}�U�UId�T�juۅ`���?�{�C�t(�į�L���R�B'�?x���޿�7P��w�vM[����7*��j8|����?�Vh��"�J�k+��!C�A���?p��ԝ���6y���O��p&X�:�C�/������2Ium�u�>�̤���w�o{ۛp��E�j�h��AV���5g���ZTVk��\퍩����߷��l[�z�T���r1�(��i���]����њVW`E�t�W^թ�&5��4���h`�����C|�g(7���]�m��I���aq�j:���d�.v�6j����H�Le%Bܴ�j��nch'�g��k+�M��o��V���s�]跊��TV!�ʹ����v ���V�1!�k�*m�*�+����.���V0tǶ�:�t^tVU������UA馲���>���\e1�fZva�Y$n��v������:���G�x]uJF���IMs�]�(E�f*������G�"�n��U�t�͜4�k�M����H0"�TV-x�"q�ʪ��M�f�`l*	��o �q�M���p�Ⱥ�s�ZxȊ���-�l������4(IM���飘Mw���H�oO_�|Z����4[[��횵�����l6�9��[�5îh�Nz�;,xև~k��Cw=x����Gw��<�����rx�.t�C�2hi0��5�6H��7g�%��*%A%�ģ�tA��t����%��JF�{�_��P0�ܻ�d��wAɘk�A�E%c��E%c��E%}�䢒>irQ�o�\T�r����L��o��y��-Wq�]�E*���ѿ|��_�>T���M� CG��oJ'�������?�<>%TXB�Ӝ�SB�ia��v��`x4�'Y����X�~�xj�����Q83��OJE�N�&H&���N� �T㘴�a��s�d��'P�]�>���K޻0&G��cpK����
��[��o Qp�1�%'_��7{�ܒ�/|Q��&{�cW�pz�eӄN.��yQ=��pKc�·�T��<��<�H���RQ�F��q��[�"
?Q=��pK]D��x��f��r�[(|��������%>H� ��?hf�(�<~��+���%_���3|�%�^�6��b
�����c>�La��v�W�g<6�WKn����_en�ۋ�����FS����<�KܞdՌ���)���w�����;�����)==e�N��){w�NO�w���)ww�MO��S~r
�Su��:���{}�T!p��j�5S���J`���	L��J��V�^+0Uܫ�z��z�S��{�ȩ^䃝L�"��"�z��z�S��{�ȩ^�^�T/�^/r�y�9Ջ�׋��E��EM������zQ�zQS���h�u���Kz����œ�fs�__\nn��y�:��/o��m���;A�J�wH؋�ͷ�����wr��z�ǰ�_�~���~o���?'�$���n��R����Lm�Z�Lzyn��"�I�?�$g��I����4�hk[��l���T^����Ƥq��n0���ƛ��Vpv���݆�v'�������&I	;����o���M{���U]��3����Osvw���&�B�t9�\�{2�,1S�^���D̔D|3T���۷���A��p��U���6?���U��[1����l��Mz�
���ٳ������׿~��W��mnƷW�d������?|v��$��e.oc:yo����4����M������x��7��w��m��ۛxs�i�G��n�C��C�2�{��`��է�L{u�l���zo����]��K����U�~�it��":�Z+���M7���7�1�{�����ft��1�?�M�������_�x�}����z�x�uu�4�mR���*WW��M�+2���'%�c'���x��xܯh<��:���f#Ւ�ܻ�}��A�l/C��ʉ:�NW�<k�ֵ�Z=�nK̦`R��H�`6R�����f�̰�忮��c�F�К:*��j�	U�T~�����FE�	���j�f��X�[�%��F>�h>��������f%?4ܓB�&�xh���G-�c�8Õ���p�m�P%�|r��4���{������7c��]�p���X�ъ�?f���ڼ�_���8�ݏ��w����S�c���������&ޜ|֟|��ۃ|�O(� ��9�E����s#����2����i\T%t��d�&�z��ֵ&pѬȱ�b���Luφu-FqXv�3�����>6f�P�:3y��b�E�x�|fD8k�s#������+n�v"[����ɾ�9��Di@m��M@/��q�<�����w��om��yG$E�"ʌx&����lϵ�5���}�Zޚ�@h�śp����^��fuR�3���S�Y��<wN���	��ʠm�T��ʻ��T�)ĲV�N��%�[R�j����%\s��y�rT���Sc�򏧜��ݬh��R��:՚ٜ��Q���`$r�5�i��~���Cm?�+�c��oK��~���ۏ�<��})�g�C�ݖ(l)��|������,�%�����0���ݘ�ߵ��Bh,D�yug6��R��FA���`*E�kKLE�����#_㟜S���<����7��f��Yێ2�.kwF��2�pjt���?w�-�ԇ7����5�E9]���-qf���`��h�I�w�Br��xE���@����,8�3��� �F�|��ԟ3�r�U��-?��d�we���a�4w\>�tZ>�n���w�ǽx<���q��~�<���#�;[��R�.f�L43[j���RS�͖�K,;�Ξ1��ԋ׸�kv-1{�Q���E��9�O���z��r�0fz��}r�ܙ��V,�zf�8�o�>�/�xs��׃�����ק�����קg_�n��Hu��}���a���'�u�w�6������7���������Ov����Ӿ�*�b��ו��U"������k���^烗�����>]�tkQ5����:��=\��՛��'k��*V�� �v�N�N��O�IΫ�U�����c�礓��}�cM��zs�=�l���|嬩V��h��H{a]nO77����ī'R���7��6�����d� �GB=#��׷�)Ħ��U�ڹ�*��L�gEt�i�tꮞ��M��b���a�'}���~���� �������˫pu=\���_����W�7���&��ޝ��δ��\��:��ɾ��4"���'�
:O��}��J�:���E��%���D��46
��ԩ
M�;%��k��9K���EU��M�L���.5A��m�E��D�FW�Ҧ64��|�W*�l{e�F��6���L������?�m�|oN^����y��N����檽|�œ��ūO�_��ޡ��?��S�����X>��~sO������O/������߾<IN�$�=y���/_onO��n7�^�˓��x�v{��:�nsy�9����Uw{���~�ݞ���Z}�=y�IË��>?~���>�?���~�Jf����Fw/�ى�|÷W�6�;������2�nS��2�3��`w�4�z�nO^�6�K,�c?gړ�m<����7���>xr����7�eof�^����<)�����?l�-�X�?���'w�%�}���͝m�?������K��}���{�}��o7W/���ɡ۝���6��Mr!��_��b�Pe'CM�^}�*��8�5쾤m��~���ƫT�ŮAO�	'N��������f.��R$"����6���O+����c���M����8��]�v�'���7�~���}�\�4f��kӿرnn��~���^�w�O�tW��K^���p������^��S���G�?�u��Y޻���؆�g��N9wE���&=Oɉ}��8����|pW��M~���Rg�������_�����
�����.�3��'�ґ�?�)�xS*��<"����Ƕ��,.��K�������,��jj�����ߘz��ٞܛ���/~~wt��^]���:�ʤ���p�ڷ����������������!����;\���e��v�������nb�H��	I����x��uIg��'<�[<�!Im������쫓6������<�m�����K���E����Ԥ��'��I�R���'��I��이�'���:���ԧ�R84��!���!�ɽC:R�?^�f:I��^nw�н������1�0������w�_&[�n�u�ýu�_ߜ���n�����'/����Y�zץ�&a�2̔��x��97r�xx��v�[�+1W�q�b�~���[=5�#�TI!����:��w�͇W��n6�8i�ݣp�C>�"|�8"8g'�5����{w���qY�S� �$ঐ@/
($0�UxJ��.���僄n��f.�z���e�����9{�<t���D�D�^r?���o"*9�<}�v��/�a�U��zwT���Q�oWwG����\�w���!�����)�|J-�ҏ�aw(�.~'`�k�7	Ԧ��١u�����_l����b�= C��F}/-}�iK����	����:�qI�z�ճ{�'��,T����`��ɬό��Sk�p����y-�����Ume^ �
��uݚ�%�EI�K��zQ��J9�z�`]h{_3��y#�i��k��̙���+��io2��&�ƨJw���M��ҺJ7��!F��/��^�A{�����#}))υ�����Wa	�ޙذ��i���/r�J�2�N���RR� g��Dܱ���-���Oվ~��TR��d����f*mυ�./,�a�m_�O�����zXm�:���?�_�Ӿ���m�*b��Cv�W7q��鯛���67q���s~�|y}3�H���?ε���K!����g�'߽t��fD����o�_P�&yb�}s���Wa�z�s~ɑӝ|ֿ�'v/kn�ї_���O��^I-��{5��)<���-d�\_J�M�~,��å�I]�/�p�m���#Mi������6(8m�g�~����2{k-������b�e�*�o��B�ԾF;
��G���mS��+nD�����Z��ԓ��M;@�.,��Fw$tT���֘�*g�0&�`L3�k���-2��RS�s6s�RϔF��֤���-����t��y�y�JCq{�.��m�q)7[*S�)�a���ϰVXj�ϛ��B�H��$��i>�%�9�g��4;�?�Y�<�.�O�RZ͇r�?�*5'u�؋����b�؋YsZ�b �[��������܋��J���ؠ�����gP�ؠ̳J�Xʸ��7�?/,��|�7�Pe�&�F��0���fwhd�v�,>�3�f��ev���D��U��R����J]+]�{��!�{��f|㱣$BtMb�K�Q)1ߛ�甲�ѣp�o�M�P�����L�2��z��"�����d�F��T�阼:�IMG{>ө�LG�g�N]�uƥ`���~N�B��{!}Gl:��t��y�2>�1�4S�uF���+ 5���J�Ϊ�|e�lҾ7��ȷ���M��J���:̿��{UXJ���8��Roݝ|���UfX��*��gZ�
TB+��]k��p}���v��n޸�..,�d���(�	�m�Kj��&���ghq&X�|���_R���q�C.+�b`e[�X�L[�Jh`3�k�h�o����|4�/+�beN���}�I�@%4�Z�I�.�+(*�be�|�ĺY,�B%4����AT��F/�JN�[��:[��j*�
V�����|sk�7X-+%��+�QTUV�t��*+
hh�?ӾV���^�5��������vST�����Ke�X��(T�5.�L�Z��U�W��Y�)�������E���c/3,
hhͰ~��@剽�i���k>hMg)+�����}#,*�d�5�/,
�h��>�W��D{4F8?e4������`��3J-�����EA�	�g��
T������7��?�������*�h�P{�)�I2pe����N�5�bz�
ֵ�q|��dm��R0oP�yRj�TBmjM�N0��!��2~�4(7���Nr�u����jde��ˌ��.����v�Uj�C/XWƋ��$ʍi�Zc�%~gT��'��e���4Sla�UV��EU4�a�(_nP+P��.�N#S��K�`L]Xl?�%�8-5oP*jm�A�ʷ2�c4(WnP+Pq��j�T=?�؟�RX�����7��q��?�T����9���7�xɜ�QW�`'�oH�A����7()����Z�����GQ%i��[ӳ�
h�Jz�=6l��������z,��I���o�ؙV��W��l�\�ף�Y��F��Ϛ>>��;��f\l?+�r�O�LF)R�d��N_�J��?3�I>�����UXla6�?V��EsQ�оh~�<�����Ypr�Ӕ[z?\}�ȩ7�����a��ӗٜn�?6��?�������>�����D_}�M����������ټ��U	"o�qu/O����''���|}u���PK   .{�Xh��;�� �0 /   images/08e4a639-d7b6-43fd-85af-03d86c8bfac2.png̺gTS]�5�R�U��+�#Jo�;��j�j齆�{BGjh!"�$�� �};��s�1���<?NF�J�^�ּ�5����KM%��L�A ������R�
0�Ջ�~]��Wѻ
���|���l��v�~.t9�����
F޺nv�P+O[
�s;{Y[���yڧb��@�� ���|ӶQ~(�����v薼�v~�f9nIy�l�0��f̂$r?^���+��^�[�{�㣫W��T�Ҙ�>�9��"�1���4���7���s��k�X[�!�x���<:��ϴVo�b����U����A��/����ۋ���3����߃_�����`���%����-���%��iɂķ�#.�^	D!��"LY.������Z��3A1�ri����	�&1�`��w�g��{e
���kp�"���Bj��H���]ޗ������t��\2d�we*�1������ᨑ�y��ˆ���[?B�\��Oq����)��M�&��D��T#}����L{|�W2}�$k���z�\	�iKiT͈�V�o�k !��h����5ÈD�ǌ�q�ǕSË~lW�����p\�Ѕ�0d����Uq]���*�V��m9ޟ:�+C�^���'���E}�a��$��O��3�_,O{E�@	��\-QS�c��_=ur����4œ\�<��X)!?�-�V��dP��CQM4\�Ff�{� �=�xS��e\ӯ���WeJ˸�D���]�`��muݛ�H��?	�b�=�e�P��).�����@�����O�&bUz�Ie�T��_0�3���C�ÿ}R������>�H�Oo�q��t۵�X����_�9�����9�R| @J�]
���╸:o�|f��v�~��`��p� d@��6��#6���t��a�v���Ҿ\�����WpM��%W4-��F=}e���y�_��<#�/�~{S8Yu�@E	bS�~�@�zS��k�P:M���*���?p'�w��ɪ�8�7��6ڴ�E>����������I�6�3���){Tp4������ݏ@�"I˙T���,Y�Tr�K?4�?�A6ʰ^Ԅ��R��|_���;D�.*<o�h:�%^\9��[���_�J�,��P�'<���~�\���Nd��ێ؎��M-���~�5@W�E-=��{����:��[Z#�� P�疍�o��Cѡ�GpS,�#�k2.���)���+��Bc(��`f��اZ?"wV7����p�XV�����i�q17�6Q孳6T1&kaΝ9g���D�M�F��|�bd�Ht�4�%E�o�E�,lz��L��R�.F����NcQ�rὢ�3N��X��
I!�eQgM�p�nV�#/��}i=����(q;����2�v�f�i!r���Me�BN��M:���'~�Y?vK�8��֏�L���U����,P�E��"2�ʉ^`�꡹��X@��2uаɅ�S1�2µ�ª2Cr�He�R���"տ� >{�x7��a���KA���'��w�k��zJ��Ee���Q͞���T�T�)���t\z�W3���A�L�_�F��L�',��L���[�z�U��'��&�M�h�Dk��Ke�Tx?6��|�U�b�Љk���O�_�����)���D��9Gݍ*�T�Y���t?^<z�N�f_���Ċg���`\�&���X��B�l3qb����9��]bz6�]�Ij,���M6|����.���U�z¤��$_�����LLR�ìw�՗H���"����/�>�.H�������6sǦ(�'o;�O�+���Nz�Y(�>[�un��'U�BY"�q��p�w�v��ja��͠�����
6�H]"�����昜s�;r2�L+|��#���8��%�f/rP�=#�����i-�_1���b��(�2��9Dݦ!��|{<)6���Z���(�gn�n5@TBH�~�Ʀ�����l�H�Y�t*Lb�^%¶��x�6��ՓH.��Q9'��P�W�����[�)�xy�f[��G�\�F��Ĕ���k���ʨ�@���C׍A����X��Ĵ�x�ß�v+�I���i�Ϩ�����(G9Bh�Z���K�)M�2Ņخ�n�\���R���]?e`
�-�$���>k5���\�Ո��:��M܍&���9@hH8��.�_���%L
 j0�[k��9Tޏ�.>�혪m��+(5:j@i��R\��9i��^W�$�=�<t �~7��W�Z�E������Ȗ�:+���F	��ߨ���5�3E���'�|��%[&�%D�Q��b�S�ώ���Q�@^K�q^[$f���oSLN�ڴ���������`�%m���$Y����ھ��-H�f`�#h��Yr�����T���;�+	:�75P"���+3��Ϗ_�x��x�k�3�2�=�pY�z�,��m*�����B��O�U���G�_�t��溜Խ�B���|�X[�w���v���U9p<%t���m���(.�(�ƕ.Up9@([�L�B�ӈ{���dݯ`3-�=�hj�`��m�����%t3Vhfp0��&�N�IR�� �в�Kym!eϹ��
���w��~���ʧm���V�9:��}*�4|�q���-M��+�f �/�:?S�@�3b!����q��;�tWgsC􆳖n����cZ}�i�8<ީ��}2��q.��#�231n�(={7�;>"[ɢL�����~�Q?ro��e��y(ϛjQ�rM�S2�y��,�O�L^�܎\�����O��:?Y���5� ���.��%=�u�Dm�����*����#��K��k�����t'0N[��������X5X����ֽ��]
��[�J��w9UZ6AAC+k����̓��[uVJ�)�����\��p3��߆�v?��S�{-ߓ��X�|�≩e4�	?SĆ5�,n�ɭ4�"����P]��C��|��n>�,���v��2�gX^��8�$��7�oA��2�D �����+������������܍\
���l��.]��ۏ6DnV���[��4S�0]|�&�r)���	eLut�N ��S{�ػ����h�p�IG]��q��YWL�ݔ�MM|(��H���MSMl�oj_D}���om��J��|H������IW/�l�6�E�U��*��$��{WNZە��j���T,�2x��A.�S&�ɬ����qځ��g'v�cmG�U!go�\
��5�n?��P��;���,�.ۆ���5��]F�/P�]1Z��Vi>?��Z S��O}B��� i-`�*��=��D��<A;}���Ծ�7􂍛�z$�a�[2A�W)qR��o���o�ژ�>�w��Z�_ uf9aϗ�;���i�l��y�ok�����*I*�j��e&am�ė&+����dɨ���h�)o�E���ǌ��,r$`n�\*I��>��6��2~_=�DJ+Q&�-s"��Y�p��sװ���nP���l�_��Y�X|W��o`�%��1��+]EU��!��Z#.�2B
�R�"5���栽D�M*���]��g���r<ف:��ohO�DeȠN�D̞��p�d�u�4�|H�i�n��&��"Z�������=yfB�v�d�F�n����֞�>�gS��C��7|�C1�����Є}���"7v����4��Gk���v��.��.�b>[Yw$Qh�G��d�<����Ud���2f�(�@_���L�"�A��~�r�e���#w���^v��-99�t�ݚ)t5�{���C����b�$��������T�n)rI��Z��J<;���;��C��Z�]!eD�1��;�Mn'�Ƃ}��E�qEz�ż� Y��� |l���G��gVu�k_�. 
�="�u���������-g���6�T�E(�0�G���q�T��S"J�$G��4;-_�^��c�w�j/*���_�<9�3:4[ߡ�n>�3�
��h�Vx���:ɸ�H?�YDw� qs��Z��������gm��'\Z�>��a�[o ��3�Aa��Ȱ*�[^�c
���֛�M�"7��3����f�7��p�)�������߬���s鋅`1����'�~
�J\��b��p�����������Rd������>�)v���'���<��P�\���H��<�i�������ݩ��K�3��>d��t^�J�������g��S��ǘ�g�Y���:;��i�V-�S)4p*c�}bG�8j|hj*�f�8�a^Hk�� �k5�$��,�VKo?٣��d��[��,������w���_ۖ�6�$�y��E���o�^�������2t�1�Pf$ �y!���oL�Gs��WV����Gt�7ޘ��[�/��8k�s�����t�\���\D��Yi+H~ƚ���������l�������A�nL�W�X�KF\��2b�2���|��2W�t
�&=����-V��k�p��$!K�g=]��ŝ��:
�j�#D���쾏�T�SZ.i�Dmʶ���r��8C��j�Y���peWe��>��t�<�zXt"��[�����)Y|�?k7~ɸ�	�V���/���T*��v���e���~�$�ճgO�j�{��PMXlj"�fe���rZ
�����P��G@GI�+'c�#��#�:��N�u?�X��@�tW��H�i8?!m��%�5Z�S����Ӿ�ܹ5 @�zo\�6��E�t�=*�#@��{F��d����!�sg[�9X@�?�z��֍C����Ɉ3�h�6�t�-��ٍ��09(����H)7���&Y[�ǭ�r�6ֺ���T,��T��,ҸӾ,�"����:�G����s���__�x�Pj^��('��҂n����(/�>��Mm����ۺe]�>�S��=�8�ߚ�]Z��Ԥi�{n�06�8��c�>�:��x�!��9�3
#J�68�\��"��,�@_�i�1�"���J�o#°l��$�����8���l M��rp��+�9ĵ����N�~�'���=?�t��Ҵ�\ƈ�s7|���� �r�^�KFx7}:�P�`��wߵVBu���F�����(��	�J�}�#=���)�
��g����ĳ����ak��3a�}=�8m���:�q�Y��C�23A�����S�m} ��)N~��:��� ��P���lgM���5�͵�ퟹw6i��_^���|��-q�/N8���Uɣ��5CM�q�~�,x��G�/��~��p��܎�i�D#h#i#�i"��]�X��EP�q�@K�kl��`.6����o�[K֛9����Ǩ����9-�o�*\��כ��t��IE��B����$���� �i�ѭ�)7r�=�\?��ڂ>� w��Jø�W*����n_q��b[����DU96�c�8?Z�R������Hw�=.'l�d����W�Ù��秈����Meƈ�����[V�j_w^Mv$��6&��W���c���,���J�.�*�w�q��2�o�]�b�&tyG ��_��ѴtF������$֝���J�-�4�J�b�/k��^˵s���j�;�]��5�9{�y捩�Q׈�t��f�U��Fy#��8^�#��-3a��0#)L
���?v>�8��65:OD�_b����.�Q�����z��Tz �د�3������ 
�ODM�8��'1}Wn�_"+ѯ��l�m�.���q,�:�v�1gqu&M����௼ oݲ�(�J	jз��V���K;���Ew��c�3{Hʳ�K ������.cdwm͙r�x��ԥӭ4�﬐ϫ��l�G^��;x���s������AA�!�v�DS��i�'5��2���fX��+	��#*Ss�D(۪�4����+r"�s\i�8sT�cpp�U�=P	����l�ʉ��9��C�ޫ�����޳:%K6�23���#E�2R
j_�Ŗ�3���`E��q�%���^�!.�)�>Ǖ�O4t5��a�c�_�(�g���#��3�X��T�/d��N�JG&;p�����?���v�
�<,���F/�Ķ��	�=(�����Q$�:I�BQ
��\����ϘN���7�aM,c����@3�}�MQ��+�^�*��(����Ҽ��I���Cu��T�A���� ~>5�8�嶩l�9����=Q9����q�K�"l!4�qV�k��?��O� $�A }h��(���@t��-�-
 �\ ��y�����Lh�7�1���ˁX��oN(���)�f��<�A� ��N˘�ݚQ�,�н�:���Z:���Ceq�˾�k`�@6�K[f`�{r̸Mp��#o���g������q�j�O���lϝX�%4g�}o�p���o����7J?�_��u�Vl��m�l�����x�q��|~6�rjz�n����Ɲ^6N�)嚢w�ݯO��#&z����ͥ���"�w"���P�� ��WO��z9�+�[5�م�y�1��/,�f��a�iA��� C���h�,`1+Ĵ�ݙf�ۢSp�������x2�@�ɼ�Q�!�[��!!��\�[�������|<ňP�-w;�P3�D �q�����`��d�+p��ߦ��"��u��aI3�²�7H�D��9�Kp�i�J2Ȧ�{�)�h=���%�����A��#%Њ�;���Z|�\��U����bU�Ҩ��SD�ʶV� h�B 	(S���K|V9�T �V���qgv�����넓n9�@w�m���-�K�� �������á_�=f����L����9����#�r�=RB,��2?ms�2u�axf`��}���Oi��^'�ʢ��o�yZ����|R=��*��k>!}�ѻ���	��+�'v&}dE
��\R�((qR��e�DsKcA5d�����3ڃ'�ps�f�f��t �l4���r0E�}�)��^R�8~Ї���.��5'����� i�H��4�y����2�1�yM���b�O5t�_�� ���#�I�9Pݼ�OH�vV���^Ǔd�����pÀ��@0��~�:�H�@}�Qp�,*���,u+�|V_0�R9�-����Cckgu>7<�8{ZQ�ɫ�{Ӓt�v��H~
#�^��B&�fj�{&I�wr��wI����jv�O�����j[��kx�`�����r�u�-{L�af�*qV%�7h}�~�59�M���K�����͕� �F��F�_� GҐ]Pc��$hr���L$����Q*l��vO���9ť�4�S%��3�:��۫k��[T�G�s����&I�ݨ����]�4���� ���I�}n[��wK���(HG���f�P.���������G�k��iII����葁c��Pys6cj���?������ο��qk�NԥE��8�_��Y����V�ܝ�%��J��f�sz��"�8=��F���6�t�hפ:�T����%qEQ���s���0~y=�"-�w���Kt��޿ܡ���Q�Q?-%`ߣ!~ZMvN藖��d�{U�����_7*|�/�J<-5���PȆ�(�#]�����G�y'胛�#�`�Q�@b�;���;C��=ɫ�k��Ӛrce49��3E1���E��R��S��bb�|D�o�|Cz75���k�@ۈ���|�\�0���<�z��g�H��r�8z�J�))J<�&���9�j%H�$�\x�&�UA?FCS̬e�g�"�t�n��_�j��$M$a�8j6hsZ�օcr�i������@7�w���� B�����^�7���ih:H��'gaX���#J�2$>G�u���}o���~�tb��f����8m��4]5�Ĝ�nGP�,M�������s;=���޸�+u�$��5�P��E�c�%�e��9:�*�(������x�&O���b5v����6�����W�����;�ޮ��O�Z��S�L���������<Z@�[�P�|[����`����nf��~$�!��qV�Ty����p-����W	"zL�e=��b��ɑ��4�:����Bȸ��߻�5����-'�U�4w9�Ҟ��ڊ����ґ�j3�G�Vv|��a���v�Os��9ǿ�h�g��R����>\�!ZV�H&�wz���E!��r�Oy�_������R ��uU���}L3�]�	���]�6t��/#��]�_��������e�mw��{���xwI��ˆ�x�C8h�J��%��RG�Y�jP��Ψ�Ȳ6t����s�5�dS=QU"�ڒ���)�˳�fmf�j��~&b��
�ܯ0�L>-�v���z0v�&kB��X"��t ŚI1'����9�dq����dtn*�P���mDS$���de���B1	��D���$t� *���<,���梋xLa�B&w�$9��[~��k/�9��{�A�lm���F\�-�Gz�1���[P�V536��TU��Q�Q�	��xH-��\\�xv挻��9�~����ϴ������T���3��;��jg��	*�!��̎ƅ�>� ����p�����Ҩ8ύ�{*	��G����:�Z�4.�/�$�c���n����s^.s�C�o�I�8dI������,O~�:X#��gA�w:f�F,��B+�eQOxH%@jB��p�8z{D�7+%��FO��7���g�!*4��m��K��@_zY�4r�~I.��A��&K�0+)��&(�kJv�@���S�ȩ�ܪ={������V��V�|�]�u,k����f0�k;قc��ҷQ�"�P	5�c�q��B��J����˛���n̢�:���Y�)p���w�~��%�Ή�y��^��(^����Q?�{� ��ڹ�;�'�� ��
��
h���+ܿ	����N���J OAw��E
�=�C�5�7Cy�>n��'n,
�[�@�{�ج�@u�A�nfjS�B#�?CA��k���=�ga����Q�AN�x���8u6��RñD��Ӄ���j��)���$NշEt-�}���ܢt�D\K�#v�U7��<�]��V'�v[%�g(��J$S+�"�&4����7z��6�1��%t���&M�,,zNZ%����i]Sb�sT��e=ḱ�/:���m ��/4#�0U=�[�!�m"6I[�D6UIX�/����^+#�ve���z�6Z��y�4�$Ӎ�A�W��v��kX���s)��<-����@�����T����9E��J�r-�&z+�5�Q!��w�8иS��\�$�����ǿ�����P�K�X�F��ܨ pK�ǐ ÌI�'kn0�a1Ċ[G,k�^cP1�_�*�o�E	l�D�EL�>9�M�Y:��g���dW~��/����f��e)۰�J�<��*��7�+Z�N��Z�@�D�b��R�}t��2j�\��>�j��T�Î�kgV����V�[����dAp�I�a�p����~��B*p�-��M DJ��u �	t��|  �r+%��^=2�N]��[+���Hz��2��s9�f��ݢ��οA�4�����q>�va��LjC{��'�8��x\M���v�ĝ ����=Hl�V5��l8�6�
��JDs���b�����N#Sk��I#�&:,��d���ޕup�?����Q�Ll�����}����������*��Pz�v��<q��f�Ǔ���Y��F�0(4��3y��6;�k����]�`�Z��d�"�_g?\kAB���ԡ&��,qFG4���H)�+�$�o��-��%�ZM�xڑ�R���g�g�7Vn���{إ�J�.KQ���{��X�IW76���M%n���g�ꄔ����LS�N�N�cS�Qc���7F:�\��P>�uFR`ǄO+�N�6�����/�=xk��z���!��Y�
"�� ����gaA驫/>F�����r�gԟ[����$����&N�ɞLŹ5D6[)�YB�2�%7��<�vj]51�u�e+G������P��;��M�����a�$�.�0Rڴ�>e���9ʧ��9"q(��Y:������V��8�\�#>*=�x���"�Za�O7��ؘ㊁i�#�Szs�o�V�E�YH<�ͿR&���$��� To�����Z�o	�������j]6��ȉz3������n�(���#<k�d���J|��!��qFh��J��XsÍ6��tL�B�U}�x9�����~�v���� ��H-bsv����kq�E�M�YE��U��B
]֠�ڂEz~Aa���@�D�������B<}��\�^4�ɠ��Y�l*���)p|�TS��R���7����hߘ�ޒ�;�ՏҨ7�i�S��t����o�pA��^rlI.������%��p�|L?�$yq���S��Wy���JY���/!$�G&\��`��?����x�6��S*�K�	�%/��!�,����BȰ�~�#�c,�l��0��y��0���y�����g,K�"�eȔ�d��h״F��?�굡q�S�a�~f�On�]�������M	�V��b!��^b�3��U��&��3��8�a����5f�~kG��tS��-���A�Q<c�D�����ѸW��P�m��E9�����`���n;�u�-T�^\㡈ɏ�V~�uC�<�]��$̧0�m3G�#	�FO���ұwi�P��IAۚ���t*L��h�o�r3�-T�<�|���#�Љ��`�O}��z��|9�=��=T�-������h��q0b�7ᩆ ����ص��W���[��IB�ͦ&�.^�5B����k��S�=���Q�~�u��J��>?��	��a٬�s�¯�3�����P>$��8��|$�<}kܻ�[�4�?��<�oI\�I5�����D��=� %�v�s}��j��*�1����Bf"5�m���N���BPo��s����*��4�:;�*��\#�ˢ�<�y�ը�#��F�y/]���FP(��ĮP
��7]���דe��U	G�w�8'�4��G3kW�s��Xe2�c�d�:��)[�p�r���㊫��<�pY��a���ΰ&�8_�o�TƔh�����wo�����ު2�ґ �0FP[t�W&���Đ������i�\�;�o0B]��/7|�F_F�ϓ볭.�����ᖎc_¦<3��)� [v�'��l���eg�����?x��u�ߤ&��d;�B�2 6ӯ�\� ��Fb�L��G�n���	�IGk���^4X�p�\��Z��vx�j��tA3�RNQ:`�F�Ψ��dg���Ty���	�,�!�U��~�W�Е���#��k��.����9��]w��1~{ŏ�äl��{N�o]Wҕ%TW�<�/����y��@C·MC~�AG�(sp�xg4�����J�� _��|�jֲ�mm�����s�7�@��T�<	"e	���()	��~�n��"Æ�f�\O�Yb���n��,�rS�� '�~��%�A=�J��M��3�Cp�b��R�#?�`u���v��ڌַ�s�n�.
��e�`|I'ƀ�����ڌ����;޿Y�~�Zq���,���۬��p��W-cnh���yYJ�VG��t�F�Ғ���َ �DJ���v����Ӳ�e{u��Ce�X�Vi�']Y�/�Y9_��c�
4=5,qV�@��4'��\������˼��N�פ:�$n��pX�;K�6ו��>�c}�"���΢��\��M����A�3O�����`�D��5�s���S�w/���Χ���Q;�Ç�T�d5u�r�rx���HS�ׅ�ۚ٩|ݦD��[0�2i�WHձ4p�1�{���U�Ѳ�3U�ǁ0���v����a����1=P~2>=���:�6:y���E��ߏ�u$�H̾zJ�r>#l���n39�)ɑ��Yn,·r���V6���e��yc�62���Rz�l�`��Os����-�r�[�)��k%�'��(ȘW	�Q�7����ٔ�a��8nDУ�8������R�v����è���Zb�'5{�P]�q癒a�_����}|���HR�/��o[t��7�ni�ĺ<);,G�>e�Y��5C-�xT���p�� 9����i�o1�S�Yxx	"t����ih��UM:#��/%����ͧߋ<��� �}2�rk��ǣH3�lΆ���)o�J۔�=R��1v`�c�˝�yt�up�d��ʷ�L��ίT�ώI~|��<BP�iذ]]Hl�o�D3}�^��`�w9U��儦��滝E�ØZglc�3��7���&W5��,�r���xC�������矵1~���K^��7�j���"��`�y�7x#!�?Nf5^_Q+�6�n��h���ȯ�zB���_�-���8�}��lf|Z�e9Lt���(#�ş�4H�Ϣ���3���x�EΪ�_S�v��L��0ϯ�t�j�'v%�z�N)�
��OD�����U���.�������Eݟ9 ��	}�8?k����	ap�KC�2LG�⾭͛c��������} �?���<9�	*z��x�I`q,�yu�����W����4��F��5��#,:�h��$f��=��o��gCwWŎ��l�X�4�v�A�F����_N�+��6e�/������D�}0�/���aLR�%|�3ջ`x�~�"S��qP�u%��đG��?darZ�Ń���:�;ˌ6���v�S�ڼ��5jG���n���g�harg���.�?/]?`}�m�3�I'Q���+Ð�e(��ʺ�d����T*|�z��2+��5l�fLr(Rzc�n�5�ݾ�R�/�[1)'qػ�������9�ã�-?�E�cp�y�\J�<g��( o9��*/4N'���y�����;�u�u���x|�k�!�=�3F*I
�w���2�Y�g����<a�B R���v�����wN^��n*^|�γ8Q�>�"m��/����/�8-u��P��4�-Hq�\��|��uA^�d����xy��B끂�}�RԆ�u�+C}�F�sW�����y�f��Gn��d���-q�����S��م,��L��-��&9����v��x�뽖��ĉ�>��Ӑ
N�u�v�IF.����jM�΄�zi��շ�.Lۧ�Q���,6ON{�56��q-��hWi~��%�Ylvpj8���$z�fr���s!P��c����Y=���^N��yU��ò7ŏҚ����L�)��k�+�����C
������*��%Ɩ��OY���KiU�-�x�kY*꣋��h҇��R<a~�>���&��j�{��t�^���!�c�Ɖ�u%��/բMQ�QW���I�[Lsf�-o}n3����o�P��=y .��6��y<�y$�A�����r`�y;|�&V����}IB��ց��e� ��/0S(X�^��g�q�OF�H�WP��c�ß�� ��
Ywg�g\�R�9��}�ו��A3UO�w%�dT ��?r#&�̆�\Ӂ��:�3a����m�����'��s��S�<dq���Wa&��N�
�W��~�ooTu����9������\����5�PÜ�[��W�����i����8`��K��0�MN�h�[4ڼ��b��}�=��lٓ�y�E���*�9J蹰�VՕ������23-����T*JF�;��B�����h�cT�NF]���M�M&gu2�¿����?nI��.�@�'>f�ӧa�u
���W񔜮h����V�����G�8>��5/���ϋ�;K=��D3��E}���2�2����W�_��� <F�y��!�CiF�S�>,��[�Q�(���k�p�Ѭ����>G:&?�����6��
n&
I��a���#�j0�<:��%���(��Rm$\{��|�v^d����o]���QiN.��a9��bi3�r����m��'X#75)"�.����_�N�9/H��:�Ap�P��\�B�d�X��?b�}��9�^z'�ҠJ�.J+�s�c�6��~O��Sg��e�)kp��ꇎ�-Y��=�z�5X�Y��X�rM�n�#T�:��X� �d�<5Yh���C�Ѩ�tX���O�֬qst�UX�)6@� O�-�+'������}��Q����0��EO���&�M&,����8j�U=��^�	D6�������(x��zN��U�r�͝�=�pނ��� ��*�*�8�?�}n쿔ε��,B|B3N�e8�)�TS�� Ƅj���=�{	�h�n8Y��e��`��V� ����u�. �M:F(O����x���<�L?�G��t�������5�핇��,#�*d�@{`�<Sp��T8^�Lm9�6x�\&r#f�@��Zp�k@|�{]�?*�%ο?�^�4�lW�'i�^�����U�\�a�O���6ØI#�s���E�-+��ק�\4�ځTT�r �Գ�PT3����l�cգǸ��n��>��_���,�G�]r=�*�yi����C���i�L[҇��t�J�����];빓�7�7�J�р��W�],NZ�͠��S��6���'R����m�t������V3�$�UP��U7��D6�R.�ק��<�D<&;��<.�d�J��n
'⬣=�%|Nˆ�|W.�!M����W=����V�=���^�'��T�+���5�\��n�����ȫ>Nf�1A�t��J⺲i2{]�:o�/{?ĸkT��(�q���8��+���]���9� �����u?+t%�x6�)����u�`�6�p413�^�n�b'w���'�r��h<3� �����s�8�]��R�Nk�=nn*v�Z��K�Ycc���mg��5'���ߢ���CϬm[��@IJA��:��p�'��Y헉���ޜW������&��8�iX ����q^ih?oiO�n��(��T����Hݻ�O�Ý.�"�7�n��_�|����p�X!�lwj��E>�k�X��L��t�/W�3���m�y�ؔ�t���)S��r�H��~�Q���i�F>=�)c����&ᥜ�#������#��S�	���m��[1VL�������WW�T�񚴨k��U���hb��`|'u�!L�x���J7SB}~-�h1I�������}�g_��=gI
R2�7�]r�C����֦{��M���O�f�_�7����N4��<�p�U�ě�;Τ;�-W+��<H�u�1z酆�7�������2�9�R/zN�f�DsE/-�UJ�b�f�L��f'�F���x��pdI��	]���yci�&�6L����l��C��#�]Ҷ�ń�1�R
#6��Fw���.���j��ޤ}�l��Yp�)]p�5�eSu�����`V�K�%�4��eT�����E���^dB[ߑ�Y�����<`Q��&:�p�@�
����.�����_`2�9,��<ߗ�`�V75�=�PԞV�_���e����JBb����w�� �B���8`3���W�7m�Vq�~���,@� N�Rײ6���ո��zS��e2*!K⶘=��C�.�ZE�R+���U`��ş�3��e �(*Z�����eυ�&?��e�i%�[Z��#��͞ɔ.y��R��j�yhX�6�a�{u����?�����Y�)����o]ux��7��9H�v��&F�^*�s���,��d*�����	��˵�$�w~�F�K{xQ����,��,E7C|�$��@�d���_u��k;�n�*�Q�Y�[���;�1�Niul�V2f��L���8����5�=}���?��*N+
�C�Ŋ�$�r�������'�[�&��y6�T�Ըֳ�25�^U������/�r�kW#���K�>6a��Uk����PDL:4��P-��W���δk�ז����ڊ�&,C��VT@0h�?���y�b�e���v&%���j�A��.܇7�.�r4���6�!8��j��!RԢ�;|�q�5�]a���%�u]�疵9��ZF��"�����T��CZ����3{V���;q>��g��s�0���3K~�kO���U��rt�a*���a��K�mq�ʨβ<��Ң/���=����Ơ`���W�-���o�ԃ5���=�޵���$��"+�4U�5�[o�R�L��~��-�.=��l�XT`�%QW��B�<���E�䤤#�tŵFm�ӑ�Pڟ:bT�a�ކ�Di�K���Žf��[|��T�����L�Մ x_}�i�k���n̝����1W���]�K�_�\�`t�5�*$�m5����S\e�S����匝*X�������d���J�ګﭓ�Cݭ{?$�O��3�SsGW�H����y�`�\$�i^����n�]��]
+PŗYt�����żWirl��i���{\��#���|;��bf�N�eT6���)EV�b�w�_-b�?=)�������\����D�3��,��nuP�# ����z^E�1E0��)���?m��߅�.>K�CͬU��g�,I|�R���1� ${=���0<�Tܟͷ�����(��õS�e�_o|!�;;�5�[0�ܺ�����?�Fb!U���2#����=����L��~�!��mM�[/�>��3T�);�'����\�Sz>����T�'��T�Ֆ]R:uߖ-�,Ȇ���U%q�j���#%�L�Gj{`��vꕜ�3Ŧ����b��|?.$}�U������O�qJ��T�)��=n+sH՚�3�ѱC��Q�������������{?~eN4?�5�fduN��C�:��D;L�ʚm'O���a���� j�{��
)�V�ݽ��V���ݡ��P��ݽh����Kp������d&���s��s��}&�ةHZ� m5˾6��m�$�t� ��R���'QƸ<���߮�z���27�-�k���0��� ��q�b����Y�LV�����_	ɉ2Q1��?����������	����|��7�����j�\����x	�kc��O�	�jMl�<�0��L���n��^�iD�Te�!�\1N�;�����_N�{�H�K�Ja�z\	�oi�.V�p�9��&y�%�Ia�s�� rv��q97;���4mI�/S�[BJ�i������D�(2��(Z�l'iw�E(�w�8=O8��������0b�sF��I���Y�6a!%�����T���
�Q<�ҏ��M%)��c=��">�����]�f{Y�Vg���iWW+����!=Z�Q�VWɏըU�aW�?P<Ib�<��JG��V��UfU���z��8�_ѧɂ%<���g���F�� s
[G��	&���c�PE�p��G ����pE���^r�Bt�J����-ͽ)��ճ���`��r<U}ŧn茴eA�)��K�_(p��/<�|�x �ېQ��b��0��"A�#*5[��շ�"3�X�`9$8}�h
A1�d5�5�_dd]X��q�n�sYo�o�:����.>�J�����o؄���(���)�b8_+ׂ׏n阬5 ǜ)����rS5Z�}B�NtqO���i�k���K��1�?�E:� �a�U�Q5#�O�v�<q�F��C&���B��Eג�JVj�+� f���	/�y�0 MM�rJ:W�)K�̷ߒ����He�~Z��ֶ/��sN�����cK`���:��ҏ��! $��Aĺ���V�ކ�Vru�7R[��N&�1T _RrfE$L0�ͱu��~���� �����Ç[���X��.ų�	\�ҩ0#1�¾��0��'�o=���'��9���[y���~=ykGPB����yؓȿߪ���4�:^WXm&�6�Ç����+�\� #޺�a\H���;��vc����}���>�R٪p��a}Z���v�<������!�8���S�ۨ����*0g�i���;"��3�'�7'����u��A�[<�5:����o����OI����E�+�:��O-��8-s���#���9o�c:���պ٬uM.m�Xj��HF��Z��4=)X:��3��ɵ1bvCw���O�� �b�z���U�����ǁ���q�vn�[n������.m=lC���8�0�m�9����]O�O���L~� a��lQԱTk���!i^$�_)��m������K�;<w����;�B��p�ۯ*o��1��m���(��emx���6!E�ɝ�������|�i���ݶ�atC_
�37�Jx�,d�D�o�ʝ=(j����]���F������Ot"zG��6z�ת�8��P�Dӎ��1����'���U��)��&8~
l���MC�,ju�3Y�������?%�_�����ܣ�����:�����i/0V�9�rsU^��۩ں^w��%����O����|\8��#���,���MA�e���o��[�҂��M`�ۚ^����-�J���L�A~7Iw=@1�ȿ��_*�ϩ��
^����uZ�<o���W*�QGl�}G�Jj��i��@z��QB����׾���',�&�dU�N�`�7�ܑ�k�lYs?��m$sv���1��n/���@១�{gc�MR����]��� �HV8� ���*Nƾ����fUi��B�L��LT��"�+iY��δ���I��PAw��s�=z�CdB1Cp������~�T�٢=oы~|������ku�2 ��s?�<2�kbE�����y��i=0��X�W���$�]�N'6~�#����R�/,v ȸ⿠��a��*�d�n���x@e��m\�lP:ة.3Š�n��/��R�\� �ۚ�'1:�V��K
8���pA��@
G�� BJ��e���^�Y�k4i���1�J�>,HČ���f��1F��J��=�ȱb�s�&D����,��po�GHe<MPH����������p��z`��{��*X]Xl�r��[�~3n�j�M�鳠���*?��ʷ��0'���/��w��wu&T��q��[�lr��1۲Z����;�,�J')���VN�(�(�Kq�z�\�:,�ٔ��`ɵ@�Ϣ�U������r�B(g.M�O�@�Ǝ��%�(P��dz=`�Cժ��B�jZ��Dђ5Ū�9�ll̓8y������a_�m�D	 5<��];�9V����ݹ�i���)0FT��E�,H�����/SNҦ���ڠS�)�]q�#{D�v��3��� *��.�u��6���ɘsH���E�X@~W�Q�r/�P)(����=j���D���Z����B�f=hC4!�z��g�Gs"r5t��:ܽ�m���+�
rD[��R��Y}�Ɓ��Ф�H��͉]��C��j��n	�iy��9��̮DG��2 �	p6��ς��<|�E-��Èe���P�q������+�Wl�|c�iB�WHmŇv���Ź�WxȂ�e����;U�`���h���k|��\ �;���e��^�,O�e�ц�K�����.�W�֛��ڗ��4E�~�L������� ���Yl�g��O�o���_x�!�.˲�:��kL���K�+en4��=>�8$|��n�n�@׼��X�5%��07]b�\i�W����r�}T�n�����N�V���$M���q?f �S��(�r�6� �q�S1uE��\��a�U�L�73}*j���f��ܡ�D��]�YQ}��ۣ�m}y�B5Aw�ZI��u?m}�OH�ܭ�0{k�q��&,���\���Zd�Pat</�m��s�7:/�h*�h:��V��11���r'���ش+��ᷧ�If���ߤ�!�}�.��������]	,�cpOd�h�ۧ��~�b�Xl���H����}&� k�>1r��Q��;�0W�,�����?�I�s)�!�5&q�Y:lk,�ݑ;)e����H;O�Y'�S�n_���~�l
��'��V���־�諺��X%��B��9�FU�$i�L����~�:�z���僘�̳��/#�l8Y����9�b[gۓ��~��B�W��g(�wg+?�v�y�T��4�@��ץJ��f����yaRE��|!=n�T�USh��oM���=�X�� 6�W;S����#^?6���Ȼ,hsW,B�D�XǊ 2g�|��T�� �(ֻk~��t��\�;`�%�/nw^�B�+� �U��ʉ�t�G~��k�r2�p��P��4!�o�j�y`�dHg�݇HG"����҃#�Ka��ސ�����xSl��,y-�>PܟH�bv�����o���{�dQ��#X)u��Z�O��F}�����閵.�Y����?��}�=�S�uyz��~_m�/��v=ҷ����ңT�z����sc���FfM�"h���I\����G��4�޸�?n�^rU?J̚�P������u��	JX�l�>��$�ն�n�����֍�j<9��IT�w��1�D�̃̔~�0>�t�,`L>�f
�#0j�� }Ѵ��D�����_ぺ��e�N�q�w�
!�4�)Q�+B���oWc#Y��hn�xB�@g�<z&��7�J��R#�542C��a�+(��tk�5k��kj�7�x�����-�ʍ�vY�aê���,x�����K���iƹ��6�O*YJT�RxV�8�M��e�MR��\�V���G9�!���ngo��2BG��d�$�?N�٤߇����|J��*�u��L��3%(�j�`�I������b��oK�s^�_��Wf0a��K����IY<�M^Rx���/���U�3~9�U'���߅��W4��L�(Ͼ���_����P�z�p0F��([��I��2�ǫ���d3��a?�܇�5������ɪV6���P��8UN�j	x#�Kؗ�DE��F���g�4��.��D�A��w���D��z��K.k8Z���B�)`�]�]�Q�arϺD���f�5�!�+��uZ���6�-��}���6�t2'x1$8i"-{��>�?}\|)y��ts�;�&<��zV.X��.x�:q��q!^��~=�ə.)�~�]�P�a��\�ÿ���,���0�_��b�<[J��_�ƿ�Q�U��'�tsjlƜb���ne�݆{��3����P��do�L͸:'���&���pPQ+�f�ǿ�<����Q�EP�1}�*����U�~f�x'W�Jeh��ΠvX$��uuZ�����2b(��D��hؽ:��"����������Be^&^<��8��Cr��NN�	�R5 \@�BA���X�M�q�p�"vaF t��Z�a�v@�(qpy�?v{!r����2�K��B! !���z+d(rn-sFd��yx��(-�m{��@
Y�d���!Y]=�ZHn� ?��@�0E��tiq�\e�y��c�jޢYh���Jb��7:�w�"M���H@ݎ�u(�z4מ0���ś	N9%�#����j�Rx%�NʠI�����+�/�DM}
2�4��c��� �"a����.:�8X���<�$��������z�8s#�P���7��\�׵5��OT��h�>���=bV���� m��on@�ceY�P���$1[���,
t����CWˁ;��^�/jS���	��-ؠdHՇɢ�m���P�����3�`Jʥ��`�a"%���b�9���ڟm����TS����f���7�s�BU���oC�����m%�¡{�k6����2�;�Ã�\��0Y�Ih�p}���,S��ѭ�0is�s$d���~�V��I�o#+v��!+N����l�n)�%ۏ����vx͆��IH��W��Z�#�fl ��
j��'��?��G�:/�\�#��]c��QF��[)I{��4�H�q��ڧ���Y��Rfdt�̵�������V����*�֖�0�g GQ�@�K��9�|��=�  qz�Q�*�R�U�L�Wb��N�hg�L*}&����rZ��܈VG�sPZ�^�<)XiF�˿�=���N������d����s�vL���C]#�[�1�I��x�*�����d�-<<�F�>�_��֚յj�z.(�s��а�KlS+̚���W�B�Y�Q��=N�W�^�l�f��P2���3� F�iVׂ.8����E����;��	��-�/鞢��4y?��5zʹ�z�T\�5���}n�̓�����q���~�ϯI\�ͩ�ѓ���lD{	:�.�g�,eL�����M��H�o����(rҖ�x}9�y�ؙ$S,�ϵ�C�����u���Ԇtu����v����N���ҝ�y>�3�d��8/}*7�Dj{���2-h��ɀ�[�{T���S!U�2�>皟�;����6ܠڐ��]��Z�� �{���<Su#�ռ(#:��N�����.YW[���N���V� H�e�נ��[mԺ�ǡ��P~`�2��&��2E]8�V�I��1N�}t,�)�}�*�8�PB�榗����ĭ���U�-�(v����;�Nze�li����r���g՞��Q:d�aY���o�km�W8�,D�yn��W�<�~�F�u�l���*���+%�	]�7��w����/F{������n^����8u�����/��I<&߭ۗ0~�|x��9������bָ�������z�J>=���{�{e�ƴ�=�-D[�+��"���N	E��_�w].q��2g�ƚ6�jiv�5֦Rl\ /�mI2WA�нi���5��������/���3���
�!�q0�il�K�A��ʈ��,ʀ�/�a^��E��|>�Խ�&�g$��ϊx�ED4!�-�߲��N�8���!�`+Q�K���\����������-}��(�l=��|�����O����u�@����@Y�����>�閜��wm�e�^��S�F�X6��ҋ8�Dʌ�
�bP�U�Z:��^h�hR��h����fՔ�സ��p�c���`��Dv�}_W?\Hb=O�+r�S��/�؅��+���n������4�8���TL���\����Fe������Ch �Ӊus~2o�q᫆��>x��H/������weI-~��J�T����:2"a�7�ND=E:��8���a����>X����<�T0�h����6���]:H��W��7
������_e�D�����THC�̫qe���aC��ڥr1�S�53�>�$rŝ��	X��(�����"��Qb,a�����Rx7W%�5}x�_���8������׹~�����{���|�ԭ��@�q`�X؈T	O�U����P��P�p�������!�B+���\����������?�GP���R6�ӏ�? ,��������7� c��o���V�.��b�t����T��˝)��C��q͹�=����Sc#E+�G_rX��������ǿ�4�H�W�3����!x��e�I�=�o�M� ���.N7�NγS���
���zM�tA�?���W���;y;Ĳ�Q��ǴGlk��jP j�ƨ񑤰�ib���N{{V�� 7�ߠ~���'�dӚIbׯ�QCĵ��m��/�k��zN<��2�V�mVI���'!�R'U�)�7�!�;���6N��V�������f�������*�j����|�FU�*ױ��M�����fċ���Ym��y]Z�D���S�ŀ�q(��F�h��2)���vI3aP�_���-��'�E3�Ծ$�IOn��n��J~�󦅓S�!>~��i�ߨ�z;t��;����������4b��Q���+�/]
�F��3�̳N���3n�X���{�d��1��"bL/���%A���e81�}��|�Y{F\Kp�6���ULG$?��U����	��v�"+r���i�Ww+=�Bd,��4���<��� �+�> �i��R����Ϯ��s��H��NXx��%��n͜�"�#/V��.=�`7c���3����Uz1L�O�LøO]�g#t���+O�Ʉ��$��g�@KzH��L�����iHl�����Q�T��U�h܃���O�r����m�aFl��M�����R���Y��qU��.
x$�ڞ��4�mT��z\��Qw�k�69���1O��%���vJ�����[�'N|d����'�XE��	�g��~��(�~֗T�V�״8����s���^����΅�,����[7&|�9Im$�i92����i�����a��q6��b(�B���+q2g:d6V�\7Һx����|�޷�#d���K�����4(��U>�,WhZoh��8���r�s�`ƻ��!lة�<E6b.T�coKsFR�J4��.Y�VC�V� A�E%d��ߝ�YKf�ذQ����2v@�{��%.l�U��'F�p���]��x?�f�C�XuuE[ye?��F?^��e��^l�F��p��|�:}���w\�*i�j��㴵��D��gʺ����Z�uL����S�E�_�prh��������ذ�FP��-鲫4ڎKM�~ԃ��j��F[���������R �,̀���{���n�
 r�g��_����LC'�u���ٶQ:�W���_ۏsT��E�!��/���e�������c� )�|��S!0h	$Ў��h>Ȧ�r��F-���\��I_�.�E��b��*��ܱtr���Rk��J7B\� �N�����Z��JՓ2�	���`X�^��M�uU��y��iW�TW��>%���5ƅO��P�)�t�������;_��+� �Q�FSK�|���U{a� ���R���p;�o�l��V�� �������݄�*)ml>l�^\P]�6���/\f��p��Q�e��q���D,�i������z,e��r��x�;�yw�&q�e��x���	Y�	�-�ߋ���A�����sv��7Hy��6�4���!�Z�r�P�E��$�<��b���<������p��oԍ�V������^��v������\-C�,@�w��������t� ���tW��?�e�"lc���\�9��ܢ�O��)�F���m�e�OL���!�LI��D�w�G�?��ܭ��vl�ɺD�ƣ�N���R'�G;�#y%B��Ԅ�r/� ;E�'��zTx�h���m�r��4�g ��o�������\�_~j���_~C�R���������2N�VoD�>�X;�!�nR~Ps��.��VY��͐��|�̜��1@}�M_Ay|ѡ7=K�K�C����|�P���H��9�G}��,!Q&]���P~Z��(;�L�����+�yxo��9��{�N�w&�$�A(�
���F�O�m�zB���lK��F���+��Cܕ�n1ǌHGxwO~ϭD��V�d����[^��%���hd۩\9RLQ��:�>�k?*
�Xa������w}����)2W6W�b�`��R�C�{��������).lb��Y�����p'5a�5���g`�,�F�a5M�Q���>��(��D{��[�'ǩ�_�#ɦ�X<C����Ro�8"���3L 4u?$�v��@�h֛<˸K>��0�:ڛભ	��� �
_�l�9��o�v��������޼�`@��)�?����֎$խ�#o���ZK���R���e�/��o��0�j��i��(I���M�v�P�_�u5V\Oz@�}�򪳚��-�V(u�j�H�KE�^�!q؈,�:� �{^Ծɤ"��y�h�5K�	�Iڭ	���z|3�s�R�]�L�
m�B��NT���k4k�M�0<���cfXQ��FŻ�t�H���'�߅�b�@�jܥ>�񶿿�8[JFk��%Q�?L�v�&����/�ٕiCW]�J7R
��bV�+��(�9*�
R�E�0�ߟTi�kq�Q�9�u�"ס[c�����i��K���HQED+��4
P���0����	�W�i���j+
�	2�R�(����f܎̙�5���+;ʐ{��W&�K��y��gocZ:?��v?�{l��Z���,�� J_����յ��8�06}�O�����W��r6����IZ����&*\��&	����4��I��LkK�{{�����`ή�F�p���:ѩ��}�t���qF,V�> �wx���2��Cd#��,9,�hϺ�_�w{Bs����搶��IkM�'�(s�D��ji��@��O��Pw�5=��*�ap��2��CO���Ϩ�*��#_B$��fI�,v�f�܏��F���� V� '��u�g�-�Ɠ������T�����F��O��+䟔���{6�ŵ�Z5�KCڊ�a�ƨQ���µ` ����*�����=u�n[������M���S5�m1��%�x�9+GΤG�}�\�邼��"i�� Lr��;��D�  $����A�W~�+oh��I^�ǲ���B�+�Yh{� ~��G968V��r�>|$w2���/
RU<t�m�[i8��	�lx,9������O����T�vf��s������t��y��[n��1�c5xd��Ͷ=��{߾,�fĘj2l�˰
�s�f���.���Hb]�7H j����&�ӌ蟀����uN[	�����zW����ML�[Cw=�>���!Ħ���������U��b�c��R���)�������!��S%b�-9�Ȝ{'�����"Z5*���B����T�Eڝc��K������\H�ω�>�T�Uⱔ_%l�;y^��Z��8�Z�N���_�E����aM �-pat����,<*W�����X>���i�b?Uk��P�°:�p�floޙUE�c_N/��u:.QX"l�̂"P�K4M}A�O�bo�P����m�~[ߏ�ڊ�0�_{�M�ᚵՉ[�(�9/֐R6�����F��a���Ň�/S�j"�S������x'���D�EN� bBPi/)�{ϰLK4�"s�ئ�`T�W�+z	#-M��S&R&�ɌQ냷	�
n�j`G�Oa��I��� ���J��cOW!*I��RIʵ��ϠI�Ⓦ�t�TϞ�ȅ@�k��`��iW�'�{��<擰Z�bΙ�Z�!�|�e��j����ȏ�Ƀ�#�Y�Px��r�`���i�$�5X��i��fƠ��/��I�z��:o8>!��Z70eq��T���^ҭ�!B�wP� ���I�������}?}��S��0�3�+DI���ͣ�FD�@�D��?�~"OH�����M5����R7N�,�9�Y8�A�`[�x�R�?!m9�uR�0�ݑ?S~\��#7�q��� ���\�,ذ��w0��:ߣ��l��0�cH!ϣW�LK�L��DV��o��x��e�h%�v�^Y)�j�W�i��������AP��x��7��{��u�"�߃�٬�"��6 Tn3J.���M�>zE�ru��8�ꯁA�KF��G�lf�4Ą�!2"���]=���`3�&֍'-T/o��S��pƚb��B��Q�|:f;��PG�izӷ��@�����ҷ^�I�'�Ŏ��>|�Gg\�v����H�$�۴���b[��(�N8
"S ��A�h%A���,嗒����W���Q"�D���ؓl�!I��T�=k~�JV�q��/75�E���R}�c�1r�̙UT5��Fop@	�K'g2Ŭ��� %��q�P���xh��	a����n��q�y��!�1�G�K�ڥ�\� �5�~��"	������U����E%l�n4}��~�m �#ЃW�m�L���aY��j�n<���:�`H��9���Q�ݼ?pH1H)���t��b���϶M��3���ƯN�t����cݢK��8lTc|��0>�z���uwi�?ވ�>�C���<7��Dd�]��/�,G�æ�0cQs�;���^��	���Y�sƠ��[+e��͸m8l0n�|���9�!	?��W�-Ʈ�~!�;Z���P��׬T:���( ����/�����VV ��x�WX Z*Z0�}9+ۃ{>뽟����e?���A�{$Vq�:"��R�9	b֠Q��K�)� ��;Q���a�ī��@��V�������DڊR�Q�hGd]Y�B1��G�bh;z��b�إa���\ߖ��͝Z��R��J�F���įq�(�:�A���;������������F����&������>!��P�	�3�r�w5����w�nDseO�-����.�@L�U}4�;�7��	y�A��� ��H���XT�2i�56�t�]0�~�o녚ւ3��cL�K�H������!k�`��C���7��L�t5pN�)Г��YK9�:&�^M�=�8B?��<�3%"��m
�x��ʢu{Ӏ$���-9�f�[a�@��[������2ܶ��*����	�7{�S�č��|�C����qԯ�p,���¼�N����(-S#N���� ޽���l��������?H�Pq�}��k/�Um-뤜|���)�^�������B�(��4��q��_؍��/N���l2�h� ]j�_{,��p�]��	(��������HY]���5wL�����~�����Y�zϾ���2�AO�R�Tݠ�ru\�J��
��	m�r��0h�m@�=��]�qZʭ]�_MC�h7ƻ[�W�ky%�.�po��*��g�H��'���iC�П,D�����;�x>i.�I{*���	�"m�Υ�->�*���K�^��j��L�4j/�jt�Y̹�/��)��l����?	_z�[.W�����_�Ux�B���KC �m6gy"�"7�cl8B�՟�������������3м�7���.�|���i�$��w$�ϫ��-Y��c��=5wf��ac�t��fAA)dz�?�������X��z�ӡʧ�"����`ת��6-zolVq�v|��*7G��=���n�ަ��IK����ǽ�_��6)��3|`����Ò���4���tQ���Г�+��~��),��XxO����B����ΘS,��rC%�H`��r�-��8�V�]Z;�c#��}�~���!�[Q/vхXl�y?�xÝ�7Bů�>��CZ@!��E����<���@M�`���>@�]���!_Et�����E��e���5]������jw��o/3-�`O�����0����
�mZ+��^ż?��V}f�7��hʓW1VT�wc�0���j�9���@�MѺrc�U�iǏ<r,��u�8�e	��5�V�Xʯ)Һ^NـQ�8:]�<��o�m���v;�.���Tqѽ�>���S�XM"Fh,�!�����@.<Vu'L��P��'Dw���gE׳j� �'��C,IM�'Y���{������9;�����Ž*��>Lm"��~���,:�2w5UZ�=��{wH��K�)�k�m�d����kge�d�����0�|�@�q�0��A%wVJ�
���jċ�Rv<�~OS�H��a5�ͧMۺ�����ۨ�!0h#���'�_�пoPΥ�[� ��G��EAR+\�5�C�������1)�-�hW�Pp�JV\��N����x�yE��g���	���/9����zL���\�>��������?*�}�r�
b���uv��	�����Q��%����>됮���T)�_��L��O�Aoь�w�|�o� F<�*��QwF�����#��2¿}�or�L�/h���5M�+]�t�Z=,�3�Ib`��qLV:��<����ӛ��S��{櫅� E���zݖ�M���v�+�w~sYR�`��=���}���5��{��6j��F�V"d5����8W2);s���WKJp#��:݋w[�m�̳z���)��^z��<���V�1��(��[��j���K�(�	e� U8�`�7i�^�^��m6{��Oy�{�BW���b��ʹ�2�^7t��%�Ѐ,h�p�Q0�p��7XY���7�e��g��WW�3j���պ�3e4i+���c7x���I�ر��Σy�|=�ms-�`�����K��=�`�|!��ˋ��|R���j�lr�x��Ꮿ@R��n-J�G�q�VKQ�xD/��z��������k�;�l�I���	aX���b����.���!�Ӵ�5�g5�!��χX�U��0�@�㞝�z����YR���n�T|q4Nn�b�p�1�s&U��l�W���������������2����aE;\��k�D>��sn!����2���ads�X8`N����iE�%�8�����Ck�~)|xΖ�N�JZi��qU�Z�����G�^�N��!��>�&���a�S��rt�������	�7�`#U+m�Ε�����ZLh���nZ�9՟uy'�&@;D�{�\���k��X�4w��7C�q��{�v���%���~1Y6j�M�8O���\o����[���[�luI�~��k��9�-a��iLD��5Ά�ԜT�rf� ����o���,��wф/���I�
�S=���H;���߰��S �EnyR�4H1A�UǾ�` �k����b�׎�%��X9 Fcg�e�;e��,oS��
�C�T5쯌N_����k��/�cn`�ڼ�F&RW�eg'���Ǯ���ӎ�*���u)*�6��ʳ;�k�� 0��z�����zg��2�����!mn�,�v���*`ޓu@��i�^�a	w��P- �͖�w`([���MO���ge��iZ5$��V�q@����Ui���j�{"�V''���xk��Ex��c�׍H0Q����	%��u܃����(��<��&�L�a�VwI�A��P�R�i��L�5D����n�"=~��Y�P�7l���X����R���WR
�7�e�������Ϸ����؅\w؆1޽$�n�u�r���ЋU��1|�Ä�Hr��Β�I{U�F��4�ma�Jȿ�$��d�cC:�f8l���Le����"�3���S�h�d�H�X�;��L����w�{�ظ�.7�2�D���|�(_K`3w�8p�r�
�]T�z5#���I	/��!'���?�՜��Ab�-��ŊxG�}�I�'��J6l�'a���o^H�<O���/�7�O����f/fR�aR{9_Ԡ��|$Qc��<�4ʂ�wS*a��55T?�#�4�F���bA����!^��̷lm'��$~�L��H�1?ܤ���D��@����Ùf��"j�5��8`2���^��	XP�s:I�(�+&�|���u�Ε�7��k����[�Х#�W��z<�����X���6FzcWɸ.ڴ�6u���G|�Dx�����5�Đ��R�F�Ǔ>��g�����^fv�Φ���&ѧdo�^�1�\���9k��A�\�ƷC�߻����i�͟��v�#zX��;琂��KW���Ut^���3�k�hv��e4���+)�t���+���~,����4�2<�˰�?}!�p���{x����aFE�~����hI@��R��OXDO8��Aڅ�Iq�󩯖��h�ֽ/-�B��P(%�e{� ŋ��i_�\|�<�gC��Co������gnj:��໥���@t�B����9�7]�!�#�
�,��@`�3P�� ���y��g��՟��C@�4d�1��!#�Rf�9"��En	-�Ԍ0��������Q�k�զ1+M��ƢɳR�B���j�	�r����k�~�17��.묾�.uw������4',kȝ�x�����9��2"�ݝx��ߌ���y�{���4�+#Hْ@I���Z��hP�n�3g1g׬Ԉ��E�ý��f\�	bE����?��� ��tk6��������rM�\�jj�V�{�����V�?d��2d&cU�T �����Q�V"&��v�\Br�&� /|¿{�npYsE�mx]VXU(�==7�}��d}�?�7\&_ㅄЈ2̮G�,s�98~?My���"�2��p�3���(�i�ԉ��	dq�&d
<>�f]���
�
A9$Rk%��W���
y�$E�XB_�W�'H��>��U�A?�@���n��o�ӎ��"�^3�F������xM���:oiG���H(ai�7^�Fq�q�
���>!�P���sb�������}�-�}�����<����'���&��J��������(��y�Kup��IBM��lXC7����\Q��?�u��Ih_QT׋$�|c�x[���������t�΁Q���BD��?�� ��<�#�E����r�͓Iw�o5�sn�-��5�Z��!��βpw-GuE�3�:]��4�0���ȰȰ�X��,����r�E�Jke;3�-�)޺;kn~��0\�g��t�����j&RĄ*���(�LKE�����Cu{����O4�mJ$���"��l�$�����Xn�)��mo��>�&�� #B�ȣ<`u��x�IU�r
��~i��m>~����$+��>�o��vx�¬�nc���b��
��b�5�BM�{4l�Ӹ*J���hc��%W�bw��[]1֗��,x�eMsZ�������8�Da���e�}V\[��+���Xr�CD��-"|*+�5G	��,E=+P�oe�G4���~�אÎC�Ā���r�H��?R7͋���Xx_�P����Q��;�;3���U�ǈ	��q7�9^�f�I���0�4�/�H\C��J���@c��Q�1>.h��
R�,
WY�Ke��g��y��P���R��s���'�9���R����m�Z��6�f����R������۫����]gB>w�+����5�g�+���������|NPx��Ǯ&@5B�����UH6� �<Q�@�O�4��j[�a�Ĉ:��������e�z.G1s]���v�PS�b�V��`��U`k����m��;�87z$/��S������Jb�&�&RnC�!�S�t��/���؅��+7�_D6�L�����}|��xG�E��!��&8�,r'13R-���鵯&�iF��=�b`Ζb}�v��v_L���1��+&#tOԶ�bNT���z���0�.���@����؊F9���c�/ƽ�R@/�炑����Wo�_!GX	f�������i�S�f|��jy/t.p�9d�. S�b���t�e���#�c
7�E�E5�$�q�vk�x����snM�<V�b�hc�ȹ�fF�r�vJ�H�G�F�IS_r���S΁���o�/����H3�范�r���g�Wo^���D�X)�|�]��c?� n�A��������ԧ�L������}貸���͝Wա2�7���z縺߸<[˶�m,�ji��Z沭�Zv-�Ɖ��9ٶ�=�s߿�����S]�O\x7P��>cpx6�8���R@�t��W�t���􅲬z��~�>V�Z����������J�
��L�'ފ9��aᕋ�ݛ��Y~�,&` Xo����&X��d�!u��a�+ځPb]+Dj�o�h߭��"RD�1���Y&h����c\���"+��D��q�R�'��L�C�5���/��j���+&P�����;�����.r�"�b�@Õ�$je<)�!�- ł�A�F2d�q�����'n��3�=~�sw�
Ne��Q�f*���Ѳ�OKÿ���uG�3�jͥ�ɠsR�5N�޴�}2���N_ 1)`��K�"���i��?I1#+ �1�G��H�_0~_M��/<M�V�g:1~L�v!����I�nU�w�ŨO�$'W�������#�~�@���5���LR\F/����7j:]O�`P*̞�:�v�|Ƴ}93}=PZ��L��������JZa�U�hHW�
&��~��2��k@U��P	�z/��h�&��� j�o"P������K���b�w��tE`dw���IS߬jܬjTb@~7F�6Q�
Q��v(H�,�_��;�1��G*�Ń.�-�x!bXA�X�B0l�9-�(6��퍄#6e93����bE ���\["v.���)^�H06�@J�X򣖛S��I�N�i����1����[��8�}:��?=��~�
��>f^ƨK��0v$��@fuP�n��r���u�'���5�~�8Xs[l	l88@�x(N�S�P�� �� ��q{-x�3��]՝��h��ŉ|�������d�҅x�KI��ᅌb�;ҝ?H�A
4�\Rq�!���ig�뵓��1ZU�����D��9�ᮬ�M��x��KA2w/t�tDK�DK�{%�!|s'��53�?\��3�J�▉�j�̙J�c�u��E���#��R$.��ڟ��.���T���x��������ٱ$pY�'��eG| �,oM]뻷
D�G��P��1R���&T��'�o eu�����a=w�g����S�;�j2����V�Z�VJo��W�9�j�7��N��:0�D"�Z�G﮵��/�J����s-��wZP fZNᆱ:�:�G�-*�:��*�U&v5U��#7{�ܩ>����t�}��gF�Q�
m	)J�F�C��@����5�j4sS+8�/�����ϰ!*�K:<��#�}.��O"m\�����8p���vgMr���~^e���EFe�!c��&Ր�j������^�����Y��V�i���)P����L���W��
^�r�(Q�a��d����f�W�k"�������q�#�e�W���/i�ٚs����PP�pQY�sY޽x�$m�:��X��g?	�$�z�0���:�ݹu��ĝ�^�/>e �Vfus"~Z��XR��ߌ<����u�^㸉xR���w�1.������a�n�R�oM3gy�[�w�#���?�8��vHC�~�I�~-]�b�}Q T_?Ve��^��q��f�@j��q����Mu�keD��	3t_�z�]s�N0���',���!�֯��V�`�_z��ebc���U�?����Y�ӑ�����QE�`-ܝ��>�s��;�܃ Dg_'�--f9�e�>/|��^����I��xJ�RT�K�[e��ѩ�e��Щ���Z/�Q�%����p��b����&���[џ�k� ���K�D3e���x�?H��G�HMw���'m97j�AY4a��p�{7jS�VR����S~��`�y���##0ӏ���.�U|>.�[��4�V���ٓ���ͩ�(#xkٞ/�λ��ʚ[�78K3�r��WM�2/���\���v䌩�V �M�z����.)�k���SJj�)�s�P���ޡb�~������J�=�A�U��^���]0u�t���3�7�b��dܒ��� ���:����2���6ˈT�u�n�i���2��x�<Bi�j��[;�EHgǍls�ٙ��l�:���`M%a;�����"�?��v�����:�X��j�#�Ò4w�HUp����։�q�"�|ÿ\��u��$�;4��i��T�a��ެ�Ǎ��p��FB�t��3҃N�H�������??r��$*W_+u�v���}�����P�����'RV�����S��p7\�y[:D������I�fj��a��Fa��1��=zYc��GL�^�7�`꼺[u�� ͅ����؍��:�Xh6y<~b���g/���Z����JT�*���٧�{�	�vn��6�&j�Г�&��o_���ML<A����n�7��$�/�h����/����P�	�!����`����-]�gi�De;�'2Cx�/8�S��2\��Dl�^G��y#�����(���cE�X�|Oϛ=�;�Bٙ�;Φ35��;��AF�%�mT��z�#K:Ԝ*�9�!=�_�הG�j��,f�� �p��ip�z��%���rh�d��։���p M_+4�Ȣ����-��Qߖ>��O-���Q�L��?~Ez��t�z;@g��6��O ��8JI�i-Tfd"�术 �����~�<W����c��}��ږ}��#����m����t�����س�6oc�ח�'C5����z�}E�ߋuu7?��X�|�Z���7���u�9�5�ҟx,�E�18p���ʥ�O��D� �^}���뮄�g�2�H�f�)�q�A(�_�:���p%��C�(!������ߢ��}XYX�	^����ԟ��1ዒ�f���kk6ܮ�QmAl�K��(�`�q�����@0w�l��E$��{�}m,	�PT=��q�������pu��B!�&��k���~ 7Եy�9���s�w[�����&#ɋ����_ۓ:0Ďj���e^<Qfѫ�	k�	2�X�Ge�k�SА�����tfu��^΂*v��QX]@1�U�����)}׍�}�re��w)�s�"�p= �b��?�<�����O�]�x/g0t��^��qҢ�{�) y8G�>>�\�@Z �i����^�@Eٌ(�!}�O=r0B�[&�Ay(���M�qG!�j�xH��B�4h,��aaqQ5i��ܴE��U��1������*L�1�S�>��=ќ8|�u��'eM�8���ך�+,���M�5���e߅a�B�� ·�C�j�I�h�E�����'�F���')#\���ד<�냞�i��)��I���8lP���2�  ��L��t#ò*����~"o�?�(���~�b�\��ox:,��j��tF<�F�;��X�e��VA9b�F���G�����C۳����(����?1!�t�K6�{���tY����PA��vG��I����<�VG���W�q.�eҦ�y/�O�b�+�mⴔ�&a*;��p�_��{v���'�5{6#�{��Q.$҅��&&��eF�3�r"Lu�vMa͉�R�s�ێ�&ΣЧP�1,U�yN����r���p��cn�JAҤް����1� �����\�-�W�y�����vq�E,<����v.79�gm�vt�*
��"M��ەI^�EM��.��{=�I�d���uc���^n��u?�פQ��A��i�
u}٬-�>�أ��2��8�g���x`1�fb����V|��M��b0)�C�^0\�b�@N	�����o�'��7U�O��8\Y�X`VAX@�\Ml����4݋�̧ou|��A]�͙����ۯ�����a�9'V'W	ٯ���X��^?��m� �|@�T�~��I��r+x�bEv��9���O|Y]ϡj(/dI�(��G�h����w�o�d�b2�ҕ��� ���H�a���@iW�$�s�R_��P>�A+0Еr<�|��O��r�a ���¼A�p̿���mlŷ:��U�C�� tz�R^����tⵂ��2�����p���A�B�9����f�ss�/���֔�T�`��6^D�щ���}�_�<#���%����y-�Q7�{����Y�|0v���V����G�?i/�os�
_b
�dr� ��{�M���,D<�1�	�@qg�v��pY���e/M-Ũ����BS\f;�����(�S�Q������ɍ�O.Hx�*�E�'��i�Ӵ�����.	3�֡�{A#aW��Uxh�AjNڠ�]Z��֓Inhum�I%���������~� tc�C�Rg���r���(<;>PP[�!p�Dfa�XM.�� �(�ep ��!:=7>�ŧ�3G�8�e�}������:�`v%x�u?u:��Ny�P�!j��kp�BI��0��)(��3SA��N�@��tO�mw��ʂ�I �
��Fۗ��#��7��_X�+���� �Ķ�e���>Ɠ��r����<תp�c(C��3ᦘ�eCi��K�3��{	c3rͩ4XeX�=&`��G�p18l]��#Bg�&#��/����!إ���*4(�Ȳ�H.GC���a&=;n��P��؋A�s��srF�e���]�z�jz��?����Lū�� ������T+���&{,�K��E��z����Vb�_93�)��$���+�>.����N0F@zs�2 Gύ*�s4i�Z)ړ��U!��2���Ln���wF�ҳ�-�Xx��1�KQ5�W�-��tӝ��~ou�e/�O�����;n��@ϡM[�u�1������W��g�����& <���ͱ*��rHR�e]���v�&���{���K8�:Ȱ%�&�iSg�l����; n�DE����z�ey�j���'PWW@w$�}k�Z�G��̝,Ν�23�B�f O<tC/H�<�LY4F4�
%���O��d�p�ؾ�]Ȍu����V��A����f��I����(�&-^+��x��}��T�24��C���8�FA-v�f���Fڍv���O�;�Kw�+���}���(�0<.��B_�'�0�� 2��ICٜ�4#U����щʿ����i��f�q��,��C���֦��Қ��c?%Wfh��>O[r�ᣰ�*LZ���5蠶��n��YCB��y0-d*�e�o�)����`o�x5��Mļ<�����s��_�cRQ�����M<�y�Nd�����
�~�Xw������Ў�]HC_f i+�z�H���Zj�  ��t�0i{"s̻�vx#q�D�}Y�ϱ����浓�%	Z�4�b�+'�BF���q�W^�|y��U�@I.���1UBb�Mֻ@�B�'&�� ��[�P�� ;m�2�h�pлv(�}�K#H��]c�pm�
d����~��d�Ǧ�f�EiE��7_�E)Qc�G�Ï�޿y�2��@Ƴj�q ޫ3�tM�@BT���{v`H}h�0<�������#���2)~s�y!_8�6D�nֳr�a�;5�M�4r���G0e�S�ɏ��*X�cy�ߗ�_��ǥغ���{����Z鼷q� ��K�g���[˘,Qx���W�J���""��$�*i���d���/���[2 F�1�*�Gw�Yu�V;�F| 8�2�5�"�g�ْ�8K��U=��&�.��.j���b�etA��Ye6�`�����>����P���� ���v��h��JĢ����+���E���vpp042"agǢ@����1u��x$�����3���my������T@l,Z��n�+����	`���"g)���g-4H��MД\x@޷k~��^���}���y��',��]�l�fy����B�Ub*/�Y�����|���hc�/�N�S�~k\��Y�M��f��X��8�H�36sͩ�'J���u�+n>�ly���
+Eq?[���v�L�=3�����֙}>ݸ��(v��N29?�A��mA�nB��WշfБc��A}� �\�w���yM�fគ�B
VVt~~~Y%%2}VbmNbmV.|�|�[K�6>ߊ��<�UU�.�]]��/�=!@�
��aF{���L�g/:��'�
���b����8�్���c%���wO��މ��m;���m�.��m�8X��^u�)d)���7��1�g���e[۽�a�ƫ��)o�������� ��z�0�B�� ���e��{<b/��d�p��'�2��GR&}�QÑc�毠�=���v'���f4�lC��O�C�wԅsܥ�bv��0�V�m��ƞ5���X,8Tp¥���"@ryu�3;;�357�&yxx�gb
�!Y�@�\����=��oڥ^�HHV���KNE�����ۊu������⧤Ux]�3�/�e`�.��B>kL��resw3���/!�B酤��Tt-�H��������O�;�ɶE(��H�V]����
}��j�ٽ#��ҰI#IG>�=�dV;ֈ��c�-y�vG�)�2����%�H�A������������ �W��.zpm)���|�2��������h�Q���W�o�iEm��Rr4g$h[qm�F5닺g�Ӝ7�SmѸ([cC�F��p��WWW�&�S��[��G!vMD ��(���c��D�����u|��S2��CW{d�YZ9ud�Z���R��Zl�޷�Á<�cw���(-;�-qO�qs�gw��}�k2�_���q��~>�%�L�
��s�	�h}�-���[�t����/����ck���.��{�,��[�;C�,1�+vJ����*�����oa����f=t˔]2J�V���y��O�~����˝!\���J��w[^���z�%M~K��Ri�l�����)(�IJJ���Q��~8��6\n�c��.�a̮*�
�Vě��f�LB""CC�B8����5k�����=l��1���U��ߕv޷�]�N�>�tx��NZJId�o�,���֚L��3A�p˱���ej55�� I?4����{�JC���X�&�^i��-zbԡ��e,��놵`Wdpp�dI��LYK��)���2�{����p��Pe�|rg`ݷ!��h�eЬ��E�yf�d�^�V��{~gF��T���?�Y�'b0�)������pZ�c7/�q$��U���3
��
�i��a��H#Z�c���e��ѫ��_!�o���|W4����Ĳ6G$���#���f:iQ��5-���̩3XR��|a�E�yة����i_����.�L��5��W}d��a?$��J���:��.�� 8e����C��ھ/U�i6S}5���\{Օ�J��LOS��b5�+���*"��G2���I�De)�h�`oŚ�w�l���_	999)��E���/��[JJjݲkP��E`4��jw�Hx��sji�_ `nq1\>�%��1��6dS�?�m�|����������bS��3�븗V�M���V���>���Ģ�����3���8M]dP��LΩTx�Ghݷ9���(�@��j f&�1�V1���Z)�r�@����>����b<5��� h�y���J�\��F��پĿ�S���Yr�:�9!<�r����S�ٓ{|d[���f6'����(Nw3\D�����U�2k�q�'�LTT ����Z̐�)��OG!�++GuZ�n8
��Doi&}>���0r���a�`�g�m��_�Ъx*w�K�j��'��bl/�Z��i%�=>���9��d�=1���{V'�HF`�Hʧw\��9`�l�O�?PA���V��T�|2�45|~tB�>z��Y�O!V��Y���
����幷p���U�&t?��S�=��c�Ff+,A�^��7I{=n���Ǿ(m��+��ѳ�[���^����!t��2]T�&��ՉK��d���0�������	��%�����S6Naُ<�d�P��]駡Ȗ���M����B�D%��D��%���o~Z��1*��7���}��b�D��|&���0�[����B%����8]�S���Jf5��]t;�*�^`���Gg1�: K�V�C$��<��,�ֺɍ�<���h#ϡ?0gs�	�fE�@Nd�V^�Z
�@��ڋ%݂���n���Q�=�^u��8y��]yڍ#�����b|}�^{�k��gb9����[m����|λ���F��$'(�y�Wg��}����nѸ�=�6�o�׏+;Rڌ*&.�:���b�wy5��N��&�Ax,y;$Hx�5���4�-���>#�īc�p���c�|Ӕ4�Q�Ss���O=WK����дV�m�/956�A�����Q�Δ�5L�W��"�|dO�,ѯ[�¤nu������'�D��E�*�������,�g���g�wd�dZe�E�I����H�j!*4.C�&�RV�T�;Ɩ�@������/�LR�ѷ�O�N�J��w<�s���rs�v��:�l8�M�uШ$A��m��H���-�Em+�/S꿍;��q������+:���X���#���(�q��f6'����
H��[k@���o�pl[��'�\Tn���yxLeZg1J�'���a̚������c��`ln]�@Gt�ŝ���͓5�U���`�'6����P����| n_���x�'P��mk�"�ru�����$�dC%M�I!�0��A�p}&�[Q5V|=��ͨf��&ŏ�������:�m�k"��/��$BR0����8C�G��}�7?"�4��<T����㕫�l������Y�J
Բ�khS,^B��H���Ң��͏ˬ�p�G��ק�<�c������o�xj�/_���6 a���bZ�%D�i�À7��)H,aB�&�U�K�`�HF# eC�!H��L��_t����,R`��y��'A��)��~��
�oy/,��Q���77����&t*N��S&Bt=9NFݕ(1�#���߆�w�8<.�)��
�
�L�LM�-՚i՚"�Nd�eddh�G�t_	EFE��)i,�BGW��p�#��B���hw�=���c	�����/c��F��2	�z|���={�	ԺAN1s�2�=fu2��&-�n\`H��ь&Mt�T`�{/R�e���V��s���E��(���:!�������`2͠��O�\�K���ޟ�S�[����ivOn�6�<��߾�t��M�9:�">B&��`�H��WVQ���8��o �H���m��퓭-���!y�qy�pu�ћ�/}W��Um��۶q�oc���#8S��5�!�$����]�OKS�o"��k������G�� 3����}Oە�I�xѱ�����j^������v�&��E��T44B��45g<����?��A�W��CX~�.	�@��``+�'I󖚋�t�z{'�wU>�$Ҧ����-tӰ���?�*�ƚ3�*y����q]n�)[.��}it0�7gٺ]��n7?D+���w�k��Y2�����#���x�����f�ok��Ǫ��@�����kX���]��ɊJ&��9T��uyyY�r�
F2p?i�Ÿ&��T�wڮ𠠡m����[]]�r�I`�0�������W��{nS.���pz�`<�[a�'2��4IO���pKRA�?��]ֈ�b\���3�	rЩP>tI~����%#��
q����'ݕG�vE0��W�Mm�O(�F� �� gUtu����r���A&�NC�u�q=Y�}e����
���~ő~E$�C��z�/$��H }(,
��u��6��T�E�G|S��d�j f��n�3�1}�o���_�V�JM��3s3Bwo�U*a��u��J�)k8�l����PV�`،�#�Wcw���{���� ����:��9���{3	�2�B��yC����-��TN�2ͪ��I���Ւ�S�}i�6��c�`=��؈+�~*ics��N�ز7��2���X������*A����/m;��u�'�,�Y���9_��yѠS�-\�)�?�ޗ�z��$c�F���X|>ſ�Z�p t2g�8 �CD�Zޅm���=������H���� 
�?e2e��	�`����7�;5;���N�;��8�-�9�8�$+ugB�`�W��ž:B�j?#̤�6�q��&��CXm�#D���'����x�ic�t�;t�`�Q�oU�`x�,Ŭ[��<M�������!�lڎ� �6҇_��*�F���5�s[�!1�)����b�1[�BB�����mx:q� ���BFOw&� MU���2M���zz�pWwٌ�����ť��>w������d2�k����J�ߧJ�u��5;���l�u�	�S�o��$uX��ɓ�.�?�A+F��\���/�۩; ��=�������&���	�޴�|٦J��Ȩ�Mbf��2e��?�|��oj2�����njq��T*>�1Q&g����a*��[��������@D�c�},�M��Lw�N�f�GLb��j5�H���V�| ̺�X�YϿ��H�)G�
��Ad�a[�aGa���t簅k�dа���c�h��A$3{�n����u�*�k9���P���m�Jqfpis3����e/k��)��7���Q�����0���E�����0���S(z��a.�4� �?f�1\�'!���,�����҇�vQXBD��/.ɥ��3޺��K�Fӝ)M9Z��y�i*R��GQQ�2���PT"�_#>:���ON�]i4ض�w�ׯ_����u1DJp/
�.�F\�4ߋ��(�q�����S����ҽ#�ہn��畍vh�>.�����������L���c��F�u[G6�)u̲��H����&��Bb;x��.��{0�դrZ������=41�?("�6��Á����=���"aa�S�E>4�d������A���c���Y�� �B4l%*h/�)����{�ά�X��TΥ� ��
l�|��1�/=r1���L����G*����N�{��Sވ�(�g`ɰ���{��H0��O�8)�`��!��݃0��֌�B�c2�2;;�m,����9���u����[���N�Cnoo�y���ഇ)��P���-O����[�WfL�c��
{_��
m�ib���2�(plW�:�5�� �v�(��G���~��%��~�l�d�p-i_�#NI1	�Z���$����2�� 8��Qy��Q3W���N.8�Z]�»c��Ե|��~g6�qb�#�w
�<����s�i�KIHq���XM��K��l�Awr%K��.����;�j����LD���Ā#�V���)�X6��Js(���Wx`]�����ƌ��W����&/��^X��30��L@���#:�¾*�,��<'��J\o�n�Y��Gk�����X|Ume��kꇀu���f�ǎD���v❝�� xeC�8���d����Ɲ�p/��󷈬n�w@o��Tm�l��~<?C�TwfmS0lTc��U�����Sj�{�-7<���_���1���@�ݠ�cs��Ŝ�B�o��j�*'w���J<����kDa}�I�s�M��H����-m�5�"de����ow,�� V�Xٍ�đ�"�����&��E�!�:�X����_��Gvѽ�)�Fjo�0��W*��o�* 2�]w��� �tFi^dj��R�y�6�N/�_Ǘr[�5I�F���Q71HVN0A9��w���rؠ������/y��"�p3���)#[!K�S�M���<$	`�v.{vk�Ubڒ�{Zi�����8��dM���D⃃�gE]lv�BQ��$/����D}f�m�2���8�h����8��6ҷ��u�A��	�L5�UA�`�L���@qi��U:T�e6����+g]z|�mߑk�&��@٭��[%�)>�7�� N�ud���cZ���!@��#>&����9�2b�D�A�:�U�p��D�Kd�q����r.�_H��#�?	
�-��RzO \H�˵���Z���jN��m���Nxf��6��Ed�P��O��$<k�FV��ѭ"#Q.x4V��U��\O�������qѽ�J��28�y���"��AA�2Mc�ŶC¡�C�ɹd&�o`	���õ�IV��Ft�U����f	�������>�����=~nFK?B���$���/�Is�j��$��U���#O2�.p��ŏl8ց|�+U{R�O�˽�׾"��g�`	x���X`�I(�O���*�TcP�׏y����cH:�� ��e�Z��/�W���!�⽤K��p��41�W@P�&�&�0���6Ձ��Y���m�,Ƒ�01f���%���Lݰf��{tg#��Ɍ�6�-���w-�{#�;�m�ʤ���ǈ�z�H�A�m[���=�+8��q�G<)�p��������mI��D�&����gĴ�)- k�5�4��e���R����ϗ�j�9z�9���-6�U��u�;�������c��(%���gt|}�ʃ��Y���x����@ \�ѵ��͗��}�DX�gd�ǫ,qx#�/�}ˉ�ͷOQMq[�gYᲺ�Lo����N�:H}���N��=���Qhꤹ��v�k�6z���Xn.��uʫ�Bx�2|�G�?	Wٲ��HÆ�k��������; {��Ңԭ?p5D�Qz��J�,][�N������|Xd���"�B� �(�Zg11 ���ׯ�1�XG��&�O�]����z�#��*�rA�JIⴐ=Y��{���>C����XPc�t�����c��-eja|QY��mj����`< �"�K�|��*Rs"[*W$k��
�g��ظ���;N?$믗S�-�ˍ���<99���|jE��Ź���5qY�&���Y%z�[Da��/K Q����d��� t~qo��Zu�Y^��B/�3Zmn�!+rz��
�7�5>OnBW��`+7��3�MH�%�ep^L�A��CCA䗒lib���oI��AF�mQ�B�VE�۞C�)3;G�y4�p�*�0�N�{�Wh��3�m���VS�ٯ���Hu���I;b�~�(+x7�#M�Z�V?Z��@�Ds�/��9�j�a4�v-��:��}�o�/����WO]�C�b����f
���is[[	E���G_1�yl�#l2�xA.X�`��J�����.��e�0U��Ow�!�ϱ�0Z�(��݄�h�������29�⛩�5�)���_e/g����&��dL�e7)�:�Bgі]/�b�k�%S���\�D���ix�J������8��r��][YF��S-]��#��Dز�9c�1�uZ	4	㞺��Æ��k��5�v!j�(R�y�\n*��8G,0k\�n�e�U��ؔv�b�}��.�o������L����?d��������c(��x#�>
�p��ZlB�M�R�'�t��[�W[/�����C�I���[<,���-{}�൩��Ku�(��7Î-����l�	VMLC4N�<3(�;`�ΘO;f�S$]�mН�W>�i~7Z�D�;���-Fz�������Aa�!mʡm!IG�bd��}B]/'�ۉJ��	}�_�KlV��G�J��Zq>�y����ഀC���dG�_g���c�5p��g
���_�vD������3�o'�L�����Z�G�����%T���	�������@��_V1�k�ti�5F���sHY#��~��)@j�|�f���tKۄ��
�m��c�n�ugT����p�!uO�Ϛ��&7�9��^�.��9���'��?8�Zvp-FW�(�K���{��� O�-x�Ļ��a�|΁�Ԅ
aF�}d&��]JD�?B��4�_&(q�	N���G���(��Z�g�ًtam�����.RW8�e��͖�O����l�|%#\^R�o2������Pwp^6l/�d�Yo Y@��"����T����e��D~�p�� ��<C5p2�0BD��������l��$�K0.瑣�9�q{�/�I�
��"��&Y�Ҳˋ
�i��ɐ����'���rB��Q�A���y���U0��>2�Į9��������Y���>a���]�挖6�]Y����0��L��A����O����m8��l��h�8���= �9k�&�2s�զO�U_`����̔�Y-��<~�n��݊>���O*n�-��!��������um�C�_��a�w��l��9z�P���>,�e�]�e_�= l�$�})_ƥ�x��`rE-�YQ'�o�ȳ�k|�Z�~�T�X��|0��{�^�%�HU9L]���������'��h��	�UYFFF@E�jdZZZs�ӗ!SS�u0l�$w^�/�@Wu�
������f[4+��4�@�'��u���M�>������x��`�Wc���o4�	��*%u�$��)SEꯉ}q�=�q�q�~�� 9�{�k3�y�����Id�_����zQ��l]
eؼ�)Cp��qZ�f�G|�� ӎ���q�;㱱5���?�����3Y��T�T�{ZHs���{��O��~ë*�8���T����t������\�fYmhj)�e"�fZ!��I�t�_0�N>2l��u�Y�꙽%ղ�%b1�kAh |�s� ^0���8x���4~_
�����d#�kƑZm���mn'��U���J���n;�M��R}�A#�=�r��>4�.F�7.o-ʹ�L*����kr��:!�|q������v�O.��z@I+*�E��(��f��ɒ���N�_�iy���O� �rm�)%!����侮��Z�:�P�{Uc��Y��\6�VLL�v�0ܺ������QY��OaZ��y��Yg��&�N�*�/��Pg��I��්ˤ�_����0f_m@jJ��3eYm6��
���8��@(A��mMػ�!G�U��?��^:�9��K�1Vjt����#1�e۝Z;���!Tv���]��:G[^?�B����o(n�����8�S� {����{��(o7Is��c����7�������I��B���'A����DAA��oUrR�;O,����
�����C[���	*�e k��7����EN̏���b�k���j�����
�W)m�x��o��K�n��tx��A� �9Uj���J"������s��Z���+ Q���d��a)����m�2��%��f<�:�4#��"VM��d��p7��[��~���΁*qo>>�P�#�x.sԷ�x(CiY �Sn��@�K)�U�R���@Q|�U�xfo9Ԗ��	����aDvf����|��W�ķTO�l��[�w�0�� <����S�FKm�ik}��B'��R+0�pF��AÔ?c����\��Bc�n��h�\�Y_���D���Y 5z�D*'�����m]����z9f��X����E��Z��,(��ʉ�{')����sH'L��ua�.���u*E0u����h�d$�����]�f63J��7.}��A�]]�J��8�.���������8['�������]��گ 鎀Z�s�����;Z����p��և=M"��ք�-�g�9�,�7�����lw��Iɮ_�2=��3����/�^�2b.��y(d���}�TR�h��&���T�d�
d`��1���=Q��W1���K��V������$�xv��y�6!S��~���aOE�$�7��0U!Ԧ����#���i^���/3����]CB�w����sG�I�+���Rs��yVE�r���t(��C����P������D�mC�ޥ��{�� P)�L}�$n���W��X{xY�p�UG��O�-�4�!�9�{騦�Ę=�O�Uϊ/�"d��|�s��m�7�qde�|X�>[��Кo�^lBa�J����7 (	y��Kdab#;���j"p�6��b����p��*!2~1���h>��8A���3�7���W�S�!D���z�#Ƕ���R�H��f����^��]�S����1�Y��1��67�]"����V�<�ж����*>������ �2�;[5꯵&-��bFy�z��p��f��9�Z����ܿ����ռ�O2,��?��b�U���u3l�mFt>]6���t,2�)aK����� ��x#e
�/A;u�c�P�s̦/?��g�o���.��#�ܩ�̓����:��쵧����l�U!�-Jo�V�'��܊�H�:h��	#��%Z��dӍ吐�/wk��7/�Kw����aҧ!��~����m���h��r�b��C���ャ;����F������<�4@5�`���Z0�b��Ҟ���u|?Rc܏t�T��}���1�� ��Z���-��l�kG,�K�&R�+G�·Hx�|�ý��*&?7��~h�d�����R���B��{�N��oT� �0l�auƸ%1�z���}�۠�89��!<~����0�U
�H�Is)�/�'�DBV?/��[f��kk�̃�6��TP0uȻ��lT7�q����jǴ{�%���&�l��k��(_�Y����׽���.��q�r�lS9�t�PW�w;����՘N�������=�F�|�;�Z�1�o�_�]]]��H���Y\�`a�Z2+�(���!A8qN_T��ɉ
=|]X$r�1�ɑ�����G�3��|�U\U��?*��tHw��� !ݍt�tw7Jw7l�;%���;�k�<���;?�x��s�9�7Ɯku����%��t7�2�J���=|��#�����>�g���.�ڼ�.�JW���os\=qc�x��Ht��r(�u`����EΥpRTs;j�� ����%.�<�Y7�L�}��R�.wH�{����2<I_�p�`���ŧ���]�c'?���FHI����?����Z����kw������<3,�9�(��<+�]����TV����߂���M��j �e�^
(�Q]�;�733����ٴ�o+k)x=�ܟ�鮴:Aт�d���p��=���]F�@�y�*|`�OD�ίIkT_�>S}K$���������#���pZj�d���NO~{%V�6��,/N�ލ�(S��Q7Rz�&�w���K%t8ꗟ.ZL�nhm;Z��#�҈1n8n�^�r%��=jC��lB�}�4���YD���{�Z��	Y��J>f���,�}�^3����=���`��lə�@��H(ʆ��^��V�?/ɹ�h�w�s�j��nN�ښGQ�=���{����%����f�����1����_��r��|��| sB�w�����_��Z����$�l��'�����nJ	4»�ǭK����,.ϩ����L�t����yrR��n��h���P�ʩ֣�Oz�=��gyޓ7��}��<���)8a�5��(�rgV�)2�PR����9�V��>�����vh]u�vG�ҏ�}4�4�o1->����-�I7c�Pb��������9H5��l�i��Tv���s���X}R�as�"�����ط���SW�~����%N���2���U;3��kY6�=��i�|����A��������8!��J2p1
��@�����ۋ@��u�qf=<�5D��$~��k�Z�k�I��dٻ��$�s��BL�,�3z��i&�;ެ�$��
�i{��n�W����޷��#x
�i		'7M�g=X��/:t�|0�z�jn�V'��"dY��J,�a�G3��r;������07�k�D�h��~r#��*���0���k� FФ>	9��kZu�=��?���J7��>�1r;�Zy"J��gc�*�Z���M���I�4u�0�����V�f�#���	��:���{ͭ�"a ��B�\��[��E&3�[)x�H��e� ����u�Rq�/2P���?��X�:�*P�����š�Ĕ�eigL���s���~�r�_�l3��i����Ѹtc���Eҹh��d�~훌���;-R��	��o�
&�ݗ�d�q[8��s��;'���'K=5O!nB���e-�{�b���#�+�_~S�.��ԭ��u��f|����Vѐ�Y���pj��ۮ��懽��N���9 �Ru����QM�{bԬq���r7(ƖK��rmd�-Yr9�.J�'��-�󳓛���6$���G{��h�br�'$��Ɖq}�/��`C��>��v��rR�^�Ae���و�Yϭ���P]�t����X�+��1ss��z߿���-ǖ�v\?���:S<�ϟΞ\��?��K��e9��U���l맪
3��'�E�Aq��3�MR]`���BZ�Ex�{>8�UH���续�J@Ta�uI��>R7��/"T���4Y�X̽��]���&�Y�T�U��a��P��
��?���PO���^��ЗI�t׃I+�8q���؟Cvo��Po)��W	��ݾp���[�K�nM��Z7?�t�9�V��x�7o��=�چ9-� ��~�\D	��G�xk�Hf�Zx�����-I٨T��;`�@�78�|��G���Χ0r��(e(1qUUU�S��}vc|�7�d���f��W��%��.%|Z=�6=^&O��/V�h&q�[b�9�-pg�.��^�	I��sQ��jzZ�zݒ�:ˑЬ��m�m Ok��K���~�F&VO#��8��S�z(�����ۣ���y+p%�ێ������܍X��^�9U����I�P��έ�ʱ��į��l��N��n�<�W@��(��\e@p �F����B�}����a��F�ԫ����JQ��H����[=��0���Wvqa�B7OO?�6�QZ��E�徭T���8�[U��6�����$����_�E��wH�u���+Aځ�����LJ���OI떊�qd���	�=�Ǖl�3cϏ{>VKU��F�]N�=p�R3V6��5"%���)�@�2>2{>2k��;BWIȂ}� !�W�l#30j���J�L����j��U�~O�;�uPj����k�X�g}D�m�����5�>��Sc�X.c�_M�mx�>�g��yv�U	T�%$��,1��Ι�����4{���7m̛Ǜ@ʳɶGR��iI���Q@�w�J��B��z�,V"o��C��2l0�E��O���F\.ݯF�NYdk�O��]�r���I�%��?�O��B��B���-��r!Q�2r��zJ�_1�}$Ff�K[�̛��vG���$�?Cy<_���E��?�qsg�� 5�pO����k~}e/t����%�4����;T�"9�`�۱ĐD�rD$�H��W���$�X1U0�-u)�v�g����I�.�:��D��8ܬ�����A��L�i��a�Ů@���c+=���sHAF�����{�J��E�=5���[�WfwF��R�`��ز{�����<�X��e<z{!IA�b� *���2O9�w((��~�j^��h�B�"�bd�$�>��Ds��@��EB	m���6����F?5q��,�Tɵ��u�/�q��6�Ƣ���~#��7�!fhkw2X̀p<N��F���btF/�����~g����+~�_�N�����AA��I߱|���E��t�����c$�( E�$	�29���nӗPw)�c�[�"��d���M��ǰ���bZ�k�`�t�NM���,x��{2��hn��~������y��$�,,�7Ӯ#�J����(b��	IƎ���5��$�!"�H�^���gA�KM�m6s�r@4]JEkٕK��q���>K)�`����z�*C,d����u�6ܥ�V�WXW�q]֣��\�SW�D���_8�?��i����El �i.}x��Ԕa�٪���YL5tt3�e��t��Z���]�(CF��ꊈǁ��v��Ov|�-q|A�'�C�d�1+,,�٨���l�Q>�Y<�#��-��s�		�Ԝ%��5L�ֆ����+q*�a��������Z�Չ[�$������I �TG@^u�)���͑P�j�H.\P��������?���j���R���������)T�re�xd����7恲>Z�e�Y��jI*4��ǂ�H�N�#{z��H�Lm�e�"��<BM��hm�pɹ�;�I:�cҊ��
+�#s�/M�>Hġ��-�X�2�-��;>\�Q*�m�ll��������!aX�v�(3b�7�X9�A��щ��k ��|}���lK����g��d��E`>��X��� =E'��Q���Ӹ�[���PN�W���f�#q^��u��PO�(���V�'��<rm=����N=T4�K��}Gj����<Q�U0�����Lv��|b����=�,cFZe���v{�yv���54$�=@׀�\�2����a˥�͈e����<��O�Srɓ�ϼ|�_��a�.�{���3�{�5����X�e�B��~��L&��0���A4�H��|>�:BJ[����c���ݗ��Y1���ga ��4�5��y����N��=��?�>RB[�tU�}�GJBrﾌ+z+h_���vP�-�/��k�m�c>F���������NQ ��O�Ks,�k��3��v"���:$,��3	����[MJ"��P�S�uq�����b�Y��S���ca�`�=v�f[�r=�zk�u���W����������2�����u������j�>��z;���KF�mػ�~~w.�LZ�j�|y����TV��xzAaa�|�Y�͆6"tt���l��?��u`��׌	:��jd�$�;�:^��=�
�����->��@�/8�eT��{{.k�Zc�n�5Λ#C�����-*��1._i9��t��"4:�WH<�C�����=��K�J��
En9f�e�����on���UT\��{�o OP��'�P�7k[�-��8�éʋ>k��W�(}��:��5 !����7%���)B�LQ���uj�����x(Q~A��bRX�Ԗ�Hu���9F�ztT�'L��힑$�e�*�wꛓ�K��4EQ�n/�IZ5�ޫ��N\�w��XQwlࣣC<i{�W�3�v� )
��aN��Y.�}#�<�6YϨ۝\��g�����>>�Ib���1z!'����$�\,�	Ѐ`�	J5C}����$��(�w��jy$.F�گOuJ�b���2����.���5�JH���懎h���v!06C�w�9ʓe��O���v�I���}�OD���sOn�Ɔ� 1���+�U{F���z�⠼)W�O.�`͞���j9l�X9��L�/\�?�:p�[BW�SҞ��5�����':Kᬐ"��c�x���1��4�FA�x>么I��6��
Fx�J�f
�����)�ML]�g�h0�7����M\ %%=�V�����IBWe���G%y��OHLL܉̶�~J����L�;�=K��>QAAA��q`p�u�a1�3]��ͬ�f�HS�����7Y�jM�;�Iint�w�X��j�#��{�<�M�	_>0,�t�7�v���緙��K}C$lDy���p���N0q�B�8����B�����R�O`�|xa�:G�E�����ڛ��K�Z��h@,�?!�{%�eJ���&�ܞ�vN��c��P�Ŋ�J+l�$��i;Wj:cxP�;T?�1���҄�ឝ��"!%�y�Ąj}c�lFݪ�Wdw�cFٰ���]2�� �T�+5��JQ]����28��'�iZ�x���+�?F3,�}GNmz�6�S�gו��W����L��ѽ�ه�L� d:?�@/t��.�W�4���n�)���P2%,�g���,jOn�|i���u�M�S��IsEb�����&���P"���JR���-%e��,ţYl�����OD7���z�`9��fh8��,���' #m���i��9�qU��Z�=ݖR� 0\��?�����b���_T1k�̔ՙ����lkk��	�)U��yG�+��.L妌�f^���kkor���e�6�3�R�
��^|P&.nH�d���jǫ�a`�� �M�#������k�XJ�ExR��������LTsJk�W�8�Lv� ��#_�Q�|T�-��pW:�U;�Dְ�c�]wY�4s'NiFo��mҿ��v�xc���bG@�
C���$�7�zv$g�B�������
eF��	��a���q�Igo���a24uu����^���8nJⲣX\Z�J��1kǁ�����Ggsjʏ&S'8� 2��͞C�kv-���}��g�]f
]T��,[z�4��,�ݹ����x�W���zg3~�K�|/�%'�YyJ��T$պ�[�`����'�E�Gh{��XJ�j�u�~��b�ܑ����/V��-��tO�L�ͭ�N#ߐ���ԃ%ǥ��ts	lq�d��_����$��b��ꅙ2�Rտ^�d�.�����q������B m�4�7M��-�;���{�K���$��,2)���etwsK��2o6�+�\�$b0�gD'W��6��?��Y����,0���MN(�u�md���dY?�����7��U;@�d�t��ٶV��%f��Ih{��W%�_ܨ�������.oUKM5�(��!Й����(�� ��y����i�P�V�]�����1�>F�jE���B���V��:`h��Q�Q��3����N//1�`���00*�\\�G/Q����~��d� ���:{���E/v��]@�L�9�:��QU��]s�>���cN���ŗ���Ϧj*��D��CT�, �~��*�J*s�\�`���1�9��Kc�1�Ќ(�K_I��c� ��~��|��������dӥFv�F� ��g��?I�l��z0e��8ɛ7o�����ؘ@����ǖ�F~3��f0�Z 	H�5��8U_6~��X�`�0�JǕ9Fnv+�ޒ\��z�^������}�>7��+¶��⬷d%��S}|j�oP͖�&��w��JJ-��B��)�l4M<�HYw��}�Y���5`�G��7������"	ko{y����f8������V?�K>#�S��q&?�i�^u2��RXZc3�_����k�ɒz�#�ƫko�F�9�)�f%�+ZEZ\!y1��OU���w�AG�1��-�%�M�������41V��k�j	�K�4��#�-G:�F����X T�`��ǒ�_���_������ް4=�,�/fLa�X�_��X���p�!Ёb&�/��S4_<]#����Uk�6��>/Yg�m�R���.�6^*페}N6��T�������c3�Vʑ�&���9/ͼ,Kr�I���AӜ\.F�%n���!v��i����:���>�)����G��$>���a�����@����?��Q\-�ߝo��U�BWoʐ��FUi<)2I�������tf�eCC=��H�yV�/P�=2��Uwo�⫲!ջ��s)8�}���fg��v�&�i��
ᷙ��qd�x��d�Q#R��4�� 2�ۇLvL�?��mO��t���EAR�������m<�����w5���/� b{}���XZ�ܧ6X�����x�����kZ،�܅����5��"�B�ZE���zS���Sj)���o5Omj���Y�L!e4�hg>�V���@t�����D�<�h���>��Dh/zd��h��Yz�O���I�D�$TP��������T:?��^��m,���>|�����%ÀG_	���,�����%1��ǃɕ�v�'1%377g�\��v9.*[(�dT��е�' GM.^-e���Шߒ�ϩ��+��8a�{a@�$��օn��s��q�E��i	���T��3��8}C��������?+p?��@l��xmA�K'����B���2XII��T���	��p$@���'�n ���c�zk���J����_��6��t���tӂS��u�A��՗��`�!oTյSr��+��̱S�ަ{��Wh~��˅>��dQ�7yLu@�Y��5i�hw���������t���w�1x����(����c4�c�&m�����p�p��I���_����t�;�+�^˫b!!!�Y�CW����0�^��dvkiR�[�p>�c�Z� rk���r	W2��S��>�&�gnHhe�!����ՒR<c xT�'�ʕC��S������qW%qSZ��b�w}�:L�Se�9��AQ�Ţ���h-�	�<Mzc��;8�ll1�,?�#]8�sň��Q��	�,P��	�\�30 ᆋ������F.���TB���"+j�����_�OM�����U(&����X�	�j5�G�g��Z�뎧L�,Dß��|��w���l�+�κYQX6G�ܧ�^�n��s��d��5�I׸��|�u;�m�5���i�֩��ii�z<p�
|�f�S�EE+������*�Ђ{���A�k;�B�NR�]Z" �PX�Q���#�ZU��E��#�����%:��ֶ3���W��z�0�׳�ŕ&7��;΅���(�=e�,�杫,t�F�4�W����C����WG�"��\�'����n��_����?a����Y/��w:�̷Ai�n�B���
�Kc���T��p>i��OA+�6���Ws�_�;������U�b`!��������/�����F�������>j���gV�l�D*�#]q\WBaL���Ҏt�7jNn3;'1�n&�V����>�}$&��X�[ݢq?f��Xk�W��LY�hc::I�z����)
��]˂��8�I���	g3�����`���f�R1c$=QùX�wz]�cɕF����"')j��\t;퀡h] ������S|��1�7�����v���Z��8n��Ku��c(-�))��e�S�������r��OVS���T���%'Ge��q�/#���l�������႗w.����!�k�5�]���-t�<�HҀ����;|��"" �/G�e�%�|d�J�N({������<��/��c^]��/�&E�n;�R���=�,[<M��Ƭ8�{:�� �����j�սo"�[�-`jZ�X� ����qp��WQK�^���rZ�:|�l6�d��l���X Y�;[.Ѕ{�d���PJ�'i�s�?�����4$:���z%k)ц=_�ǚ��ۦ�rF���������,��U���5������2����9�6n��-��h��ԟ�����BC}CCC���*T�Ui})"�6d�p�=�=&>O����!��)����>5Wd��\�Z�[�	�d�8Ek��I�)��3�%��2ͤ�A"�u~p-�n�l7N��4]�D�u�P/:��J�u��E��\̑%0���
n(����_zJ�^	 ����Y�Cj�GZZZ`����?���0ۻ�����A�i��/o���+J�W�M���������ؼ��S�oҍi%��t��9mFF���"�g)Q�U��ٱ�ö~Q����B@-�3٣ugnp� @�Rs���g��������ߞᮁ��Z��C~Kl�!�;�D������!����o
�ˏ WR����팲�"
$.j;{���yo�]�����8����*�2�BE��o�b�b�p��������JO����a���Xw�&�j����@��
�o��*�r�5��V?uY�e�N'vn��$e�S�����}q�$��[�oy�� ��lԷ7	�\g�^��w��Ο�s�Z !d���L]QL�� |"�
HXTk�ⱱ��v�:`#���9�?���$s뚓���d��ӧO���BA�qp@�>�%��2x�TB�rI�*D���������D:1R�6����0��i�-�4��j���R��>�pM��qPN��*ޅ
���"H��D���#��;���>�9��%�\!j��k(�E�a9��_T��v9���|��&KT�~���h^�x������IQ���n���Q��g,�Ʀ�O|��]w���u�����5���s3��!Y)��4nz3��x�1�h�	���z�u��3�?�r���*c�=u�CƇ��$�@>�䞤�w"�N���[���8�mv*�?���"��Ũ-H.0]w��C5�wQl[�X#���,` Z:���4�Ûm�����E��-�oB��~��a��j��,ˋ_v��Lǳ��GS����c���^������SY�g�	]|kr���̏���v󒵏�����h�_'7̪d�m�� �t0�f�j��B��ՅS1y������U�{z���B��ʢx�W`_</�h�j��,
/��߭���RGz��s�FZ�TD?�L��Yw���.9����lf�{���n"����� _.�����阛S#E&��f3t5�&{�����K��[r��Imjx�׶6Q�,���q�fѡ:����9/$o}���a=����r}�A�B}X��W�ح��x�X��22��>���&�:~F�.�y�4�� �$��cJ�4�g@�:��$pCG�J6�(�k%�s��d���@I�-}�I+�D"p�`Ee�0��|��B��t=�zsiq����a�oy��~��NnP+��ϥ}�����9����L���6Qc+'�{��BlU�u�w�{z�b����ED��a���w=i.>�4o�HBI֥�:V���n9��p���hd�v�c�d�]����`d��D<��e���/<��� �e�=��=LÿȨ` 0�b�R&�^ĴK)����T��CV����֊@�u��#��$Q�]8�޻&fp��jQ�^�˛����r�"�>�+$"�|�r�۠wH{�}0��<i�s@�s�F� [�o�"�?����سPOS4a�����w(p��)�]·��f����,����b�8���
���=���-T+Ȳz�+*P�{�>YZ��a�S�.]���!|�zp��ߙZ�П�$��c�&�^����bfF)��֣d)��!Kh�����Y�	]4;x-c)��<��
����(P�uhhi�U4�<���3,'��0=�]�Y�_R@DP����S��W��>����A�.�ЪW��,(��E~f����+������k�B�e���vJ�,;f����%��M�i�_߬���ֱ���$�BV4u�)��!��E�dP �:�3�k�[�P���0&��#'c�+� ;7 ���%�]]��J?	��8�'1S�а,e���O>P �g��u���� �Ɔq�3X}ѥ݅�ʎINN��i�o��hة�:��t�4Jk��!N�k�4�B�D�b�z��R�d�>�^���}�{��+^�R�s~hCR-�;�O�TYU�><�/pk�k������&�v%��K��C���R�[�-?�w�M[�շmxXn7�?��y�#�H��oX3����c��������vX0�����i9u��u�Ӵ�B��4�:k�:����>6�U��m5>��P��Qmu�l^�8����4���k'�c^w<'����A ���g��m��g�� tU���s"�� �jc����W�α�+�ndL⭜���m����Z:[K7M��FU9�R4��� ̊� Ê
�ៜ�<�(ъM6н�!!����?q����\��ձs��J�z>��-���p���$:`�N�΢>�6x�u��q��'���� ���w	��ʃ���.y�sOB�KIFe�7���K��i>-SH�����c� D�^���0� 뵻�h���+y-M�fU�hm�<>M��%����&OV�ؽ��%牑!���P�ִ2�H�3��
����B>��rۡ���q;w��Nd��!r��7E�2��g+K��	�Ǉ'ڰ��"ـ�@@�Ʀ�+ɀ���F��2����4�<!¾�c�6L���J�m'bm'*�ӖO��O���W�U�r�%��7�h����m��0wK����w�t��]q&�7%Gfx����<:L��DU�s" R׋��nLm�����Ʀ�qF1��(��Ș=�p��K�(r�@{6��u�6��
4t7J��]���x�'f��"b|JJ�x,Ef݌���?�?�r`�Ku�z�d3jPS}����,ܟݝ�'I8^���-z�$�*ܜW�}�u���q�y�xQ�j

��m9��Y�3&����2a8��+��v�x6u������e���+���ӽ���PV�!i˚�a�;��/=���b��z�Qyؙ�R��(s�Ġ���Z����²iũ��w.]|�"�2�fL���l��2eg�M���l�Ƈw�-+�����6p����?���K3�-,ҡ�o��t ��40 �Ÿ�gmH��!򤼵�9��_�� p�T�)Y��=�¯�����;2h5�m�e�����=����DE���s��gp$�kj��ܥJ[���۔�Y�~��<���n�P!N����/EI<6/�+$�*Q�"����X�`�da��47���Y���0Q����b�Y�q����Mg�(��f����Xv� -���`)_�]�Z���J���Z�.���ΚЪԔR��pٍ�y���������c�FD�B~���1��$,��D�a8�:l{0����Y���D5y'��if��r>���ĵ�q�p�oܷ�����0X|P!��ěz�k�f����;6����ܙ�&��N���.���E�؁ӵ@"

p�KبT�'-mW<��T}j�ܷY��/7�oDy~���MC��?U�J�H�7��i�yi}o&ט.
�X
!��,&EBhG[�r��_��OB�EΚz:0^����9�F�VE����`�k�ۑj���p8��3ty�4Ӧh�x�����m{$�jA	���p��RB��!�p��O��Q=�B�Wr3r|��E@�=����Z����S��O�x�W��nN���--�`�e��t�k<�Q�>���ӊ��K�78W�H��D�5n���b �(R]����i����E~�vDB^�}laa̵ie��1^�u���%_�l������H�+��}�/�C��A�D-^�0gs	��e�w['�PSS�'�/}>D�x����/��"\�Zi^��N@����р���W�s#>	0c�CQ|IK�W�����`��s�a��D��7�?+���Ǒ�����Gh�n��K��lawet�Τ
���1_�sr�;�rLH���#�F�M��wR"[W����	z�+�u�o�ҟ�Es�u�/�N��Y�o_Q|������.pR��O���I����b*���� �{77R�U �Ζ��p��2֡>�nM��<�s��&�`b����Ȝ;27uʦ�0d�6��
�n�����?�B�H�ʃ�s`i���h�05߰��R�b,3_-oNO�)��^��fM�J&**:����F��Sf �T���'���Cp	��HVg̒�?�� �@f��,4b���0��v�͉�w���92|�p����(�;ulP��@��䵩�}�2��РY/(R�c#b�RO��
��I�W�:�jt�͸f
���U�]^�~,b�G��S~jj����l+!�"
:�q����&��no�Ŭ�9E��Lx"���L����$	��
� ��#�\��_��"���b*�]F+3�j���%�A�9��] b��<\���Şb��¯LL��"Ѐ��l�~r��X���M.{��8����ej��7�F_Du��.e��Rv��X�-39B<���11��k�9C5v�k͵N�a�L��|�����"C�,~k�7s��gc^�C����� ����7���c :�Ń��Pz�,}���s#tkÚ{.���$��������{<5+��6����*�p{/)k�cPp����Lϗg��
�f��>�(:U11�5zy�V�D�1w,��DA������)���s����蚋VÔ]L����;��W��ױ�(K���TJ��v'��,�9_HO��(Yz���=?�Ht�j��@U�����=��p�������̌���$'?���M�eM�޼��S���xf���@�?XFq=��b����-E#P���}��r�?�p�s��O����-(p�F�Q)��ى��I��I]���ӌ���1K4��ا��yMʂ�"�"�$�K��&+x�.D��[�K|�Ncp�~f��܁Y%�#�[rz�|GW���eU�/����@ez���C�"_m_LiC�'�-d�(�����#�W	��I��8e27?�7_����$��d4�����G�H�p�=��؜���?�r"��աnN��K]�Dbuoc-�H�\S�*u����IW�d�ϼ����)� i�l@;�As:<9"�J�j���_�����o�hg�H��;��.�������å~��o{^*�Ǫ����N���]�+�a�&����?WvQ1�u�gBgma��^�����$�����ܮр�U�D����ť�͜�[�9�<�p�ʉ�21�N�8 ���B�D=]���<����k������׽���6�»W.��>�;����R��Eg^�4����y
�?�u]�L�`-��pQ���o�ُ�?�r�((C����M7��f��C�ڮ�"�Ӂ%����+Mwoo������}=z�W��M�����~܉�a�D��$����W��� ��6��qf�����,��\А��a[S#��v{�>	��e[-�'Ի��3�eG4�	K�`կa�`��N�℅��g+I�ܯu1_r7���i�YVW���G���B�@ �	�U<X�(���P�D�S��G�8f��VQ�%�[l�h��ϖ��lS"[��މVT�vH!ϯ��寿�G��N6OX��r��}}(���*0�B�1q$_H�Z3U"/��LH�bNIk`F$~��N�t�$U����bMք�`S����� �%?տO�D�·�w�=	����U�*U
�c�Ϙ<�h�w�b����[�x U�:5P���>f�v��U�^�]k�w�N��L]���8�ᗆ�|<4>�̬��bb�.Ą]��A�ǐRl���x� �p��s]y�
Ma��/>���҂���u�����ޓ 8��`�U��f��Ghf�L�����M�N��0�=�B����NI��D���D�O����Ӏ{����>W������v����z�PIs�j�,Q*��p��������ө�s/t9i��~�V����7��Bw��¡�w6�u/\V��o�E�zx)�12�h�vqÒ���-�>�"���L���uJ��%pG(�th�����X����I dꫵ�B��>�E@G�U��z2���S+�@�$�P1}����Id$�}�Mp?-���j��S��ۻL;{D�Ǝ��}���q���/}�o�ϫkҰ����.�{�cO �5�97F�Ĵ~����P �{C4��NHxG���п}�0;�O*���U�͛�v�>r5�h���I��)e*��.1Ck��'�f�҃�W+(Z]����u+-�*����z�?w��^�/<5P�����2G�c�K��6UD@�	O�^�m]WI�xԿ�7�q��\oG�w�8j���֦�N��l�!��P�0���ޱ��S��2**��n�t�U�I�"|�2e]��f?8!.��}�{ϗ��W�AS=���Kk��؀�a�xt�ohnf̺�b�͉�'DV��ǯ B�i��#�斖�"����W��ڶ����bJ�D)?���ׯU~�SY��X�NY��.�-U��a� �r�{W�>5N��P,
ԉ�'�2��v�b2�Ġeay�	�L��q�a���WI�b�&3h������s2z�y����C=--��D
��z ���������������K����jL4	g�`�[(ʋ���B�휫6�NJ���&��k��[����α)?�>@Ѐ>��fI�"$1;�2&����}��T��~���8�ri�\)���wս=@�)�/]�.������3-�N������M|Po;W�Ẽ�5NR��4+��7e�DH�b����Hf�6w�6=��)��z��˦q��wd*%�
ʦ���9�!c'*J+��R�{AKD8	����c�ᩣ/cZUh���1@~���r ��S��D!'���e
��bS(	��'��T�WB�d���#O^:�����e{����y�{��wtd�=��f�Z�(��N�Og,�(�{�)b���lǳj���A�xl�}=��|!��Lg���)H��\�%���5RG�8����*�m]���D°��	������~�=׫l� ���56��q��������+.�����f�_&(����X�ώ��#���ܛ[�Ɔ3�9P��!�^窞ܲK}nKU���p$� :�a�w�d��o� miS�})
urOA��ȶ_[���C)e9��f�+��Q�����Q�>��U)K��$��}BUs�F�e���P�:b��Lkqc)�}�o��U{w��N���Fˋ�/88*��65���H|v+�|�O<nQ�<c�7Ёb�,����R�9�:����T'�ppp�o�~��TA�RV(�����ME���%���r�vp¨Gb:���oMAi���[ ��O%�pA1��r�����x{��.�-�7B�|���>��'�6�S;����&�!3��N+3�SN̢]��`UKD�eê:}gm���X6|�DR\��S�_vmB�b�:j����dEY�=/�r�,�8�hk�����ʒc�Q�A�@GR̴^]N_��Hgo�2.}�L�zV=���!T���\�`<��R��dR/__R��[�:;�Q��� �Z-o��Qy�͢�f��xr��~Ѻ��y���L�X)�~����u- ��_R%0c�톯�k����߫�%N�6�p�U&�Ouu���*@i��Mk�_K���j|�<�����Q���&B��o*��p`F�)j��B�puu���΁9(\N���F��	' ��GTQ�gX"���O_����tA��C1o�����f`?��L-9߹�k0�~��r�/�Dh�^�*�9�j��̬��cJ�ʷ+k�L�
�'��R�$���N<=�5i9�o�b�b��\��
2�z���	�M@G�#4�=r����2�?.�fW��5k��"c��Sm���+�ĖUS�zl�yx�.�o��S��&�<T�T�<��G&�|�)�Ga�wi!���dMˊ�2$�E���NEK�ݡôG�+ǉ��|ט ��3,<����K���8��G]�v��i�*+wƙ+�A)M�x��/�X��fX"����\��Б�v�NUj=[���MS��UV���.�t~�0����;K�A�ꞈ�"F���z���%N9k$T1�e�C��S <��J`���>6�W�QW��|߭d������'pc<"e�>',�8}�'�-�c�}�?4�s��� |IX��Dh�t�C�`�_���e��SX��t�W>�����2VcC��?+�(��#��ᾦ4� �x>C���Y}���|ˌ+�PE�+:�7!s,�Y���E7m��ˌt�M5k?��my���C���v8_3���������~�e�q�0������%͢���Q�s�EUZbq���p�Q��jd�O��<s�=У�֎���ϡ�0���[N��A�j|y2����qJ3�Z�C�����Vl>����Ԏ�[_�U�u�"��H�R�Hw��"�����ݝR""��%%���]�9���{��;�y�^{���\{�}RL���<^�V�_2��k��Y0��.<�ϳ�[M������Ғ_��p��%���KeX!��6-f<K�[�,�v߿�n?T�lZ(�t�>���gu��\O�x����A);/��c`����9�h�'� �+�?�?VQ��i�(H���ڬ\��}���TVFM?�U�H���&��wx?� a��R������r�FV��NϨS��v�Gq@D������N�I!W���R���r�L
��P	�����9�J�EX�:t����bh_���Z-@틃���Y����ƈ�:j'�M+*��W=��3�>�%s�Zt]=ll��!w8/�𩘳�S�Y
��c���O�f�'�>ңK}f�g����Y[		�C�����F�1�S,�L*+�u^���A��*+�u�i�ވr���nȞ����hW^55��o%�����V}��U�WZ��-7��x{:^l�*�g~�X�fcYYY ���?e���{PFXѩo�7f�[��{�8$Wl�����9�o5|wO���DzH��I����J��4
[}VJ��]���r���C��Z��!j��=:9��\��!rw3�<_:K/�e�a|Y����M��C/��F�þR�Ӣ��WgpT��&�V�D�i2��Z�����gf3ծ���f"�]�'��$O<=a���0��i;�K�-w����#�nk(�MUb��N#��;�?NQ�p9!''_XjjA�������Jz���~�M�[��و:mWgCʼ�}A�!6�KL�H)֢��G.�lq�o��ϻ�b_+M���@�D����s���C���A�3���4�2���j|�����(<k�c7>0��=w��www����n�c�.��]f3��\����f��8?.8~�7G�����L�<<�9�Wx�+����E���� ��2(���)�����H�g��J��sp!�~���&X��L�h 4���;ȈauU��n�<ء�NU��O7�T�6�3��G��K�~�4��Д��¦�q��	xl���X�tm�L �a*D`-ͪ�DM;���=d�nLeR�������f�^�m���.+]b0Iᕺ�y��J�T�����wy���~J����E���S��;�60��H��D[P!��y#�/�F�اK	�r���nH@��쫋I����;Qh���h��K�7o��o�~*����!?�l��5��~���l����t����w�cRH
�3����v������/@L{؞_�)U;�XQPCr0dH�Ū�����tA9Yn�ؒ�"d{N��N�u}�~��fnn�����M��L��>�-����=� ���ܜTA?B�/�JJK�����J����ci��|�*�lbQ��A���O�m˝@HP���|��3���� �@��60P0���D��:$J ������t�Q�67W90�*l^��1�t���]DO��/�H�Ϩ��X��������D��ku�06�zxl��R�[��ޯ���c�T]�6������V@Ja���k6$Z�b�h���������D������n��L����LJ��#�B'(��7��}e&aؿ�y_��Y����%l4!͎y?���[  �ڢ�(��~��"ĆOS8���s�\y���C0Y�� �m'#LT!41���&�{�H������ X��l�E��UV(���U��fp
;n��\��}}�W�0Bm��c@�M��	�x�5F(�X�!E���M��</�V�Wx8Q~��	�@����Ѩ̕b��G�E&'�3��|�.`r8G�%�(2z�1?ET�Q�%�$��н�ʾq�mk�J>:�����@(��&өV�5}�)��V��+Y�QhH
�b$g�Td|ȴ�G�w�PN9f��0�)}"#�Z	r���8�b�~��)�;�%�h��K�@X�������fg˾S��:5y�1�/&��3�G ���	x� a��^�*���%���'�>��%�Dj����d��}�z���OF٣@����c<y�#�=*<D�k[[5y{[?L��=a�E�#�ɣ19?y�*u�{)���s�2��T�>��jw��k#��}�0p^�����/l������pgCD݆o�Y�9�ȗ��WW�@썡�+.������D��U� #;^�Yͷ�50�zܷ����A^]�3���ȑ���>M��5�Žŀ�^��^︰0�S���yb�u^�
�DX�%�5����'}}(=��-�����Ia�7\��fϜ���CUMu���s�=Kk�/I�\�x���x���_�i���3�r��Dqǧ��|y������������LD�cJEupj�3v����%!�q����%jc+O�������=[-�����=e+��踌�D�P&����[����g!����DC���.��}l���d�TOS뜷-�^ʇk�ܵ�%D�I�9U�e�Q�n��g�^\���,0����{��X��5�����5���[\{�}T����e8�K�G[	�xdpQ;I�[Q�����ǲ�߮o�ݶ��E���oX�ڹ C�*�� �wW����!!t��/�,=Q|Ёle�^����t��;�*��w��N�����������[X��������]�VY���I���:xu{�(\^Y�(��
��}H^�9�i}MZ�sj��8+� "V�L�ƒb�ցL��������x�/�̨�(��/&J>!������o�ް�q=�� �����`|=�PѦV"[T\	'Cg���㫕���͎9ۑ����(J��5*��y?2?�P����V���m��r�|�c�������`�6���s]������k˄#3ςEaB�8�3�P�f��|�s�wuu����/���ݼ/A�>�p���30CUCЍ�≖<�I�/�&�NG%����P8�y��ɧ���(`�~�������5�q�w}�+�����3ֺ���`T�\y�=�`nMh����߅^�v�$Ȍ��e�]0�(��£�Ϗ����ٸ��������F-�f��o�󏙆�
;t�B��9)��
^��E{��$4�(���=���)���r���	*g������4����0Z�����R�A=�78[�aFb��nS�Y����԰S�94�+;O(���d��D���]Ӝi��6��H�M7�!�&(��D�9�0dND��se���}W���|�}a��{���<SG���>F(ǆ��	������#�}����\���W�YH��_y�.O����k��v�]R��z��'ZC�4Dhb�į�PP�����7����;�2���6���;�_����F�IF�i��:<>N,���21Rfݣ+^I��M��{�;�/��w5���x�yg{��gf��� 󢊑 �/"u3B��I3�Q�X��iB�c����s�B�\Ը��i�ϲ�w���_��")�۽�s����+(�a���~�B)(��h���~�]Zc����~�yQrl�%�utr�L6u1fA�����4��#��U{8'-�x�!�R~c��X�U��-� ��?� Xԛ	�o�+5�xV���=]_83�Ѻ�?��t��e���Q�x_��L����E|ݘ�U'!��ע��V�����#�q%������E="�X�d4��$}_��;џ��~Q�CRU�P�������<� 0����t����QHG��s���p}#��(�\a[5���-���X��I1⯙�f���c���H�_�D�-�5�Oh��,��L){6���g�o��s}Xi���94�5������d�g3�ƭ��	�x�܁[��o��L�p6m����Ux�[N->q���|r��V��w��m�R����}5|fpK�
3�;�8�����bIX�T}�1
G�Ll�	՗[[����������Q��@��\�C�y��魬�ҽB��F�RPPP��hr0�x�q�����J��^��aMZ�C��~�ʫf�^��柹�T<S�A2K�7Q����Ef����B�,У�f��M�xT����jvjBmE3\\Z����8<����A�l��3�wl8������?T����,.����pt�_�����O�7qӾ~���K�R�X/�m�d~20�+7i{d5#�?S.� ���Dg֥�e�NF��J��ۮ�<������ܵV+{�橴��*Ǜ��BK���ƛ� #��x�u�����l�՗/�^Q�-
��	��ea��	�=wd������2���_|�f�C����[#ԟK�Ѽ�����(-��]��C��`ñ�B�,���N�:-
t/ 6���"���鏗Fǥ7��uf��/֔W>��g��W������u\�Y�=�u}�w?�?y�ş-�����s��N{��\��9����΄�w�.%w�ޢ�$Ll� 6Uƹ_��L�vS�}-)�[�e�G�^� n�<6��6k.i�!��1vZ�E�"m��1%S��vk����,K�#řb�J��YZٵ�|$�����CᧆWQ�[c\$���m�N�Ƌn���4M��=�]�"�
�c�1�s�.�+G|ՙ��|�+�9�?a��l�%�a"h��ak�q��t�a��ܥE
��$
�pP>�T��<ܖ8G.ײ����qW7��E���� 3�Ɖ�̛lԖ�~��rf���B�ܬ���������c����ƥ��1(-#�O�J��dͦ�{>�xwRk�NA����e:&�����w4"7���g�d�n�r�O��]3�=�꘿sFI����ǁD�/��@ 	#?>�-���|��7�����JI8Q`ѫ�~�~&��^\}ux7m�|]���v����Qu������x�D<��*u0"�R�)�&��N��K���K[�Ye�z��dTz��&�9;;�YYY_��:R�{��tr�f5:���������-J�a����7r#1��&	�G#��ɜ8y�k\��4�{<�_ ������2�0Q��W,u�{��R0C���ʰ|V�.ҠV�S�$��j�sxx<8�M�p6�#�~Q��1{�;�wwn�;4b b�qfe@�(K֮�DDEu�~*O�EeٹE�W�k]�69���F�{�hk۞�b��������y a�.++K�٠�z�r��qBB�ݾʮhQ�8z%�%����_��6د;�n��xnUi�q�\]^�N�i��j����^�L�i�Fg�}v���S�	mL[i�I�;���{AM�E�E�q��kgA�[����W~��O�w�B�V��M�,�7$�΀A|���F���e���##��{��?e_���a�xޥ�ŝ��*b��q������.�=o�S*�wU&���pb�������PF�>U�[1�sɐ�K8�ȳsZ��-�7�0���ך;���>����8n��(U�Q���6a�����r�R�Ԧ��D7����T�5�Z�XXgWd:QO!*?7ȇ{��#Y�{���23<����2r�?�-!@����J�ܿa���ۍ���9��&u�~z�.�2[a_���pwl6kgo�s����O#�js�q o���υ��#�5~����P@�F�$� Z4���| k�$7JH�C�|Wo_C�TWgqu�i��������;^�'��b�֖���~Z���=��BA�J<�GŘBTÚ{�a��
�����í�jZ'৬`8Sj-�� ���]�Z�d��J��2&>�@�)���a�c!I!pjD{�e$u �/�p(�é�LO�h�qk1��-6ǭI>����w�����ՓY��i
?��i�y��824O�u}�-�r��X&�M]9����H�y �
���s������%-L����;���	��'�y��aQ���UG�3.�)m.�D��lm۶F�[���	�&3*w���wW����lǹِlZ�v�˓����"D���od�(P�P��֒%t�\$���s���{����!\�����泽ޭ�_�ˈ�	�K&��yz����F
t]'��"J�4W�������{����i ���}��/�X-�v@]���A�����b5^���\4t��ы.��ӿ��@����c�:��
��64*���W۴j�"$@?�{� ��NOO�I�4�֨361Xݛ�^00��v�lY�A�˭�|���)Uh��O�,=��B��t�HJxH)�},$��q�=�e��B����Q�;dn��1��z���$ddD��j@LϬ'�uu�@��&�S	.�����n�m��� 7S4��q�'`�N������툧��Um��B�M$�W'�S@t�L��|@^����VTVv�h�^�h��Lvq��b�@3��c���>ԠC
	����)��<˕��<.�xf׆{�����.$
�ԇ+�vr�f8����]E�^}�J><ay�xRO�l�2{Ѓ�e_|s4�/]:'g'(γ&ޮ�&C�9v�`R�`�Jm�SS`2��(C���^�O����f��}�mC�D�5�;���T)$v�2��6��>�����2���(�U����.;�K�\�
ep?|Qe�>�x!QUSz
S��'hh�}��n���t��Bjk%*����z}��'H�=}}(+��!��+�^�QF��}��N֤��&#,�+�_)���(��T�m(������	�����"�4�9��%Tp�E�1������q�j�-/
��F'ޅ������h��s�[$�41UgS&�m������*�qgpdzÂS��®��>�����F������7��-�����&�(��0?~��ŧ��� C�֦io���P(b;�x�--����8�����٢���SƗ�<U�����8���;M��wgC���� 49:>�`a�f���;P{�է��%�����S9�+h�P�?|�s��`>!�����Gר�� 2ٖ{�-��v%^�/rϜ�L�k���r�7���n99�w

�@:!a�VMLLX:q��T��;L$�I�����V��r��gs��v�%�A�dd3� �%׏�M��ogX)#� 6��B��g��:Zߺ��>��Y"}\�!t7���@��6��|q+�Z�h�H`g��3��b��mM������l�uu�n���P=��,�-..���9�����<nj�$��D\�;v���	��~@$������5'�pZIQpq�300L4�7nP�㸤��q+�Q0[��>��SuZ7�=V���������^K W��$�w����m��<�9r{,��x�m�=�]��3�[XD���FDD�!�|�ƛ��B�P�F������J>���k!����BT<|����<�=��k��������rީ�ye~�QR!���%`��v�&~���W����!�
^�X"B����:ű����չ쉌@6`8���9f���
@/�H�����4�_UUӝ,����y�}���5��^"�A�M�+(�cI��{�Ei�Y��Ht����,H@󃣗���m�Fw�B�Y�ld� ME��$��w�f��qTS_���|�Z��ο~��;�EBE2o���7���h�� ��17���Ͽ��&��&	�^ ̔��3G����������9s�y`��0s����g����\^\�N.�3�;ڵ�V#������eG�����|dlf$����?��wxԍ�����Q@wWW��Z��wy�ncdJffL�����+ r�n��f�˥5�T�,�0j�.4�e<�r�b\x��뵱�[23�Yt%ӳ�qk���g��?a�����D���ͻ��0kWu>��  pPο��!���Û�#)q�a���Y�r�~�,A����%zAi�j�l9��)�o�ԩkZD@��ny�.�rY��	���f=n����4:�.o�Q��N�=��L��3RD*(*R���d�<�q�׼��U���T������[Z0�w�+mA�N�l[�x;-�wT�\��ܦl�_`#��R'�]ph~Bp�J��"�/�@?W)A�)����ɀ��U��d C��+RE��w@��I���9����KRVV,���O�4Tk�e;��%,L����Җ�LKv���a�_�]F��D��}��!6����x�����0�\#i�Zt�Zԅn[TK���a��iv�2�IN�H�Y'p[ 0��ǝ��&��S�o@#">�Қ�1�DHP0<&��C��X�`-��ظ�NB襧Ì�{|���#lk{�v�[�<͋��C���Nd��o벼J����9�l�6����i��� F>��\(��j�S�T"������,==(%* �c�>�zb;��y�9U� D����w���e�6�4�8�gl�Q���+�	�����x�l��fF&���������G޸ ��D0�MPb��)�]kWM�>����r��=���R��{Xs�bR}���O���V�M�+p.]'S9�ʂ��-�:��O=q�؇��y�p5 �8� N`{�,7`���3Ua1��E����e� q2���x�2/�`�
PR����m,�6����>m�5w��Q��ѓ`�r�'rnL�{W�P�$_`n..%-����)�M\�g���za?���'����J�R=K��-R��Ef�4��ao'<HW�###ш�^s�ugeW??�?�dp)$�Ѵ}�����GW�]M�׽�{q�T��:8��\�y���KLOxi��C]�;6����O���;���\r����ի�{C��u�7	S�'�y��*��cr�&�������~=θ>z��f�Gp���W=�M4?���PBC��R��4\J�4/�sҚ��/.zְ����j�T��r>����9k8R.<!�o���
S���[�l9��ȗ�{E��?����J�3A�=���j�X�]�3�������`��������Ka!���-��9�`1}�r@Ꮽ�L.Q�HB���2���p\"��c{�K�����v�`���[���y8u�&
� ʭ~��\?���i��y����^A-�g5�Uf�6D���-5��;#F˼F3# `��ܚ�	� ���(����������RKS�x�"ҕf�k��2��u.��l�S��F��i��,RZ�ܒ��W7�'���a2#�r��	o#qI1k'8SSӗ��q���˧�b�ε��H�T�g�����N5����#3�;y���(wեr���'o�����r���v�u�O��b#�1�r�M:�677�l��&~��To �x+����]��U��X�&��}gg�򂡢�i�=������c��W���N�� ���ئ����*�����'@f���M���:]����p<(27FP�g�_�7,G�Y��tx�l\R�Q�	,��,�ZX�yN6����'�Y�����6�N��R�*䵏������H�̢�=[���,��9�:v��SDj�nƵ���I�"�R~�ܿ"H\.�޸7e�'ܣ����/�"�����}rN���Q�~7{9��VB����%cI��l1rkIP��f��~N'��t��� ����]��e������q?z�K쑞����j1
(bɌ�%%�	n��+@�ު�?�6�${�E����i���Y�����5.= �zkk�Ll���_G�G%Id�eK+ �	���A���˗" 9���#��9��-�|�hS��
X�銦�~�ň���E����,,�̗���$����D��Wv�����N�'�3�Ljj������r1X�8�ӎ�W�$/�0p9�N�b�R�d�1�D� �8c���s�:'��Y�Dq�i��z�U	���@yynFt�9����_���p����H��Y�ٵ�&0\��3UcN�qT���l�	I��S�O�8�^���
�+����,�-Rk/m��p@�]�j�aw��RQ�<U	���p�
���@���?��BĤgC&/��j֧Od\����"�1����;n1A �A6���D����vOa vj�O����
��^0�8 �< 3yI�))�[k(9��f��01vځ^�
�>���1�ݹ=�h�C|�{v9�٣�����9�>ٌ����H@U��Jb��`s]�"��i������<.3�yЌ�� ˣO���D$5��jj�z�������{L���N��]�ٜ�2��k�Y��b��|�r���(��#.�a!�z;q$���!6bDZ�GpԾ�X�l��W��H�w�ߚ~{��&A!�'���ŕ%$EE6�ꪦ����g�b�*+��9���`�m�j���ت�Y���4�>����̾��,������gO�kz�θ Z/r�p8G�FBB����Fv���dLl��V�Q?([���Eגd�@z]Ã�,b�"�0����yǫb1��wC ����eiQ�ScѫSd�]��X2S�xG���ٙ�����a�����,Q�xU��C!��f�o���'&=�Ƕ�5�Bw�?���)����P�_�J��[�µNO�'���!����XX`L�Cu�V�9��o�E���	`WS*�?�Y87�%%:��, r�7��#�ϸ�5&Ό�&%�/*���\����X���:���s"YW
h���|$��4��_�0�����=�9b��8�_��}>h��d���Sɵ����R��x�|����ߛ��+,t�ޡ�}�Pl�.3����
uq�5!�ȎG��V52��9�ˋ�����sA+#�۝��M�A��&M0 ʵ�����oA@���r&rzJ�X	P+j�PӡR�[�J���B���b@���+3C4#��KL6~�hs�� ����R;���^��'N�p�ևA�e(p���FL��{�
���,�>����О��0������ͫ4';��ѣ��Q~e?i�99z䆇hU�������L�Ѥ$Vu6���(Y���j�)����v�T'���qwR�����N��|�(���5,:r�'�YZ&~i3׈uw�|��"��*��1yoL�\�}�˙Y�7e�c0��H�ep��{���3�d�� �����Я�~����r��z,����t���v�3��B��J��|o�h�e������W��L�qJ����D��RH,_��������YKl7w�$�%cSSQ�YX��12-���͍�xS��9�\��z��v�ybj
J�Jrl�i����L�.��^ =C%(4�vii	�	�<cаJ�ɂX3��hfs���������=�m�
�g&��0��󇧆��"ѕ���gg��Cw�<=2X������J���R1g�"b���?�}
���K�ّ������)i������l�Oʦ��9�*��#���SZ~�x��]sF@�&�asq��{���iY�}��:Sm�/�?�@7�y��p$�?�}zq�������NL���M�@K�,a��#���Ӥ�ќ�Oyo��v��Wspr�4�N��l_�t����W�z�#,��F�ҀV����I_0W^B!�2~��̈���h�&[�����>��@iTbN���=a��ׅA��E�ާ���KH�A0ttv�n�p�fJЁ���h:�j�Ub�5z~��M>'{�2ɹ�����6=��5����\\y"�;�۵YЍEҟ���{�S�2(3g穨���.G�[Ŧ������ ����� %Y//	{����g�&*6(�@��u��� �ݳO�\�GO�-�{��P'?���F�ihj���S!�_
lЧ?��x�J�����!�j��/����B�7}|���f�־�L�\��~����b��a-'c e �����o�b$��;H�(���n��6H�544���N����zK�-ј��%�j_�嗌�}�Fq�ڎm�{ޣ`�RT7������NX�$���l��:Eɾ���^�I"��=wJ�' ����t�N��0��M�� �~
/&6�� �GGGEF� �v��}ۯ��r�� �rj�GT�3��Vl
�%3��L����QL&�{����`��okk'c%}�p�!]N��S�/o|EO,��:cY)��G?䱖�Ic;{ۅ|����9��ע���#?|������*K��\a�2(ܗ��Qh�f�]������	,v~٢!��3��p<8;��lr�����mb��`)�����U[�<y%�.�Qj��l� ��6;;���GHx��Zh70^�W?��������/&��3[B��Ag�$�r<d���О>�%#g�������7T�ף2�p�]�����������7�I.�{꼡�w>�o�5�^��	��<N���M��葩��u��8ecD9��K�}�Pa��������U� �+/gW�y�#�RSd015�$s��h
�{�D���;8��jk[Z�1}�{У����?d-(T���LJ�V2����&"{�D��JE����^�������eD5@�����9�*�6j9�Ƿoo� ��7xp�"�ЭG� ��t@�����{5�ý����׎�<ǀ�{ q���� ���Q��=.�)�o��03gZQ�1�t@Qe��͉`ff��Y닷�\-I�[i�.���i��;��gH��ĻP�\,-����J�0�\���>Ļ��(죍�M_�ߖ��O�l��#��`��8�576�`+��H���KH��-�c�9�7����$���}Ȅ|�]2ee�@Pz2�P_��٧{��4&�� ��OM��~�P3�	�Xd>����?ڟ��&��l��Ui$���)e�A/��,M��yY�[�'�e`���d �5a���,;�*g��P���*Q��AS���F})\؅W4W������5 �_ �S���3�?<&6���y0�������{ee�Q��ӆ^�0 �T+��zF�RE>��������+%d�yyE�(*!,�ɦہ�a{tcNE'u��b�>
���rɠ�3��(kk��q͇z��'a���	���N�ſk�|`]HGUU5��B|:g;�;�����}cJɔ��/7��"�c1+܎Ch��h���g�̊�ÂD�  Q&#�����'#���J�U.�/~����Cu4<<����4���Y� j��~z~-K�vfϺ:n����S�tT}򗜉�U1�]�\�%L�D�J����I`��Q���g5K]�"�ƒ�Z塭��'J	�����?$�H7<==�B��)�::�`K�Ŝ�Qɠ�宅�2�[��w�l���x��j�_TO
Q��y�5lwo��-�\�x��Jh�j�F����SXx�����&F@��?���3��>UWGJ	e��z�xw���9����m44R7�	c,-��}d��.�b�T���s�k��s��%#�`�+�5�op-9��X��3cG�MQ�iE���2���Լ��I�Xb�ާ�A�#nn�]4� ylRby���?ןN�bZ=�3�m���Vykô��_�Yaoo�?(,�R���sr�� ��r����G���22X����v�V�,�l���� ���UH3o���ݐC�V#�,�o��.M`x�he}=�t۲ş�%C��̹�ZI�����*d	``ji/�P���!�(��#a1�ց��
]YYi��}�7����4�H�Q֡Ϸ�MWp�p������0JNA��g/	�έms V[N�Ȩ��[$P(�j��Y}}}�HD�Zȕ=H�CD��a"�<lJ�־���Ou�$�yG� X�>�(�l�r�M��X� �u��ث�s�.LLL����遟}���������=�È�����(��P��Y6*IBggg�-�>����P�yl���ظ�a���k J���
swvN΃�O`���	y����;�g�[��f��$''�嶂@?())�%����Ɠ	��y���{���7��͝	�1�oͮ�'�$�����G����#��r�&�L��� �b{�}p��ǣsk{�y�O��k,�����<�=DE��H98���ʐ<��@3���QJ#������A&����q���L	���e`A/IG-���K.'=_,���׬�X���`�@�[�������o"H@<LlsL�(ᕏ���h��>LQ~|�N�0[���ژ�XXD�Gn��a�^�>��	��x0�[jL��J�(/{���U�Y0�����[��d˸��m���.�d> ���� �5''�F�m�&+I��	���!����}�c���_�Ie�S�����777����U%;:����U)1Q^��gl'�������Z��F���Y耞+*�������'�1��M����[]��7<
��*'��%��5���!@X��Q* ����՜[2���/م�H]f�'>ufd&��Γ�R:���6�\X����a	�Oֿ��d�U�E�����>G�����޷Ύ ;�z��N���r'�d	^�y��\���S�� [c���|--��������Q�~֬�;ZT^�hb�D��v��<�<	��������'*-��-��r~�	�zDٽ���	�`y��e/��3B���	L��Y^Wɫ�C�u��N�7$�?�/�d�eT���Ȉ���Ԍ��ŉ��$�!-DEB �5�b|J1��S�r�p�ݽ�9����J�G���y>
�M�-���4 <�LW�ed�㾧~!v$��Ŷ�5������yr�>>���B�k��l������gW�K�m��	2�;�
´X�N�;�Rj̦� ��(Lo41Cy	۳��bG�m�����������R�
�ך�_"�N3t�t�9(���iF��KP�Eٔ�7M�E[���������,k���$ijՖx~`�/���-�v���BE-��/��]銘���3a.�2���s�{+i��j~aص�i~��G۾��%�[< �Gtu�����//!�Q�ܜ��hjX���C4�Ĕx'';{�333�ŕ?G����F��y��NQ=
ݛ|�]t��х�[�9CI�l���-Q)����b�1�5���]+��oK���[-�ڬBYa=: ��6��Pk5�6Ke-'oiUj��k�)noo7����[3{ۛ�*mi�p���{gu�(�_�7	�!�y��V0$99��ݦ�s���.l��?2,W�h�艊��sxr��{�qR[�����F���k��mB��Zuy�D�;����c�>�iV��y2qj)��(��D�	��p���`���i6�Z��+&!���g|ؘ�|
ͅ.#:�BT`Ŝ�������)p�W��k�~~
�;lT<�������
��c��9��������n:.�B�K�".�����Z5wM��c��W퉪�aii�z�s��&w�k���U8`;&�`�������omgC{$�ƫY�ȵ�?�to��i0//��P��ga��q����k� �+�?K��[|7��W7��FI�s^�^2�L���}s{���rJc2M^( ��	��Ȩ�rtҽ$��={Q�ݗ_	*I[�4|�;4��{��m#�ɪ���_�r)���U�x����a���8�H�n�o}�%K�s�3�ƀ�|�/,/E�l���C_�'��Skx1��3�d�ӘR�IU�d�+%~��k�,�~��.��F����� ��uߍ��J�1s,�4=PZ�~�y�Z�jd���z��3$��u�쑡�5J`�	� ތ����~�����,;}J�Ћ��\���c6�߸FaA�}'&��d)>ج�q;](>��)yM+�8�([��J���H� �n��9�qU��<:@E�V�f��a�*%#Ӷ��3O��V�׶MMP���vM)%�-p?:��ܹY%�3����;m�m������ i�:�JJ�A�.�d^;tY��79�Q�&&fFV�_����o���R,����f���ZX��|��4�5-�HMM=8<l�,5 R� ����u9��`Ⱦ�_�#_�Y��Ŧf��\#G􅖃#{H�~8ߨ���u�w�E��3ka�8�������x����\1B��(�cp����[�K�Ʈz/O��I�PN���G Ѣ�Hh��E�'(����W��i	#���6����&I�!�z���0�q1�=|�^G�O9 ۾w(�"nlD�:���$���(���y���S���m��X����b��Qrx�	6k��|>.{NX�JNK�@��'�T����2�2@��nˏ�g��h:U-:��,#�E��?�du=����,Q�õ%��v�U��D�"�����Zr�xwW��$�G'x��\s.�U�5��x%x���^V]V�����f�f���.?�!$�9Z����tR�����y˪{���³���e=+Q���b���o|kܪ}�Ŕ�z��m�Ƞ��v[�.�Q^oM�D���TD����R�ŊiZ�?j�������,�@�b����@b0`��
�vbW_��g��}`F?�~T�2z;�m��F���`Y��n�Y�i��c����l[����P��Y�����P ����UYx����֮�EMx��C��l����/xK�{^p���ʩ���kc!�h&��������/���}���(�W{�C�{�Z��e��J�F�9gxEZU�)�
s�Z�ۏ��F�)2!jν�CK��:�#�B~i�Yu�'�p�L"��5�k>i�2;���n#)�=��v�-����|L��A�K�f�����Q��^� ?]�\@���z���1���]u;���w� z�֌ْ�
R��ǹV�����o�$�p4�ѻ�����d\&��J���}��ק���!�i�+ �0�;�5@#��5��ɉ����|�O��Ds�C�#�r��741�6�{��D�����l~�(�5-�f��V�;��SBK� *N��"��ר���o�c��\N�ש覾����I��7ewƺ�y���kq��)�����4��йt��N\��o�AE184���xm���(h\e}
���gM����S��+�F���Zn�{8dptwoAw�8v���l䳛���e��텝�vaoP���5��'��oR	-���A�d~�y��_N�o0``�R4tB��;����|���E}�B���s������{k��b�l}jD�	槟�ة�o yF�_\G/F�����تI �B�b�������(�GIf_����Y�W�U���F9�F��ʒsך�Z�Ob��� �7Y��BxhX3D7��4{���r�gc���m\olj�SQ�%�v���v�G;i�O���ugq؇M�|��bb~�H��3�K�~�e�@%���!��H����uù�X ��7k0���B4�Y�SoWׄ�b�݃����I�5�� �$�CAwww�����p6��s�TQ5�W��ϻv���oa3��e�,�Ry�����+R���mj��Ӂ��a���|�i^������?R��,$�6=����W�����&z��$��a�جR4���������[x2��¾�������u�`�WĻ�2+�:@#d~��s��m����9U1�ѵt����%S���dHS�LlL�bª�d�@4.j�l-*)���PG��oz݋ɢ�@�=KG�����Yq�O�ӵ5�z%�LVk�
u��GO/���_�׳gO�ޙ�_����5�o���2�0��_�n��J�0�C�_� K}}�ͣ���qXz���z�4��`����D[���Q�6W:�8N%���-%{=��� I��/ԡ�.���w'���*�U2�G�a�kk@��C�)
#�Mnw�};�Z�P2�d1���l-{��F�	��� �I�� ���W:�����h�-Ŭ!�������C�#L��u�n�q�6�^
�*fh)+hu�i�����^�@�^]7ǉ����ᐗ�^Gy���!��c=��p/��F�D�y:���/���IB'�U�:M�+�j����)���qZ����-#�"A����U�c�Gx)�}��:SF�%�ɨ$~�
1�٦����"#soF|P�:�����CM�
J�3��v���䤥3�qA��W�k�������9%%-�7Xx�0�a�4����RZ-�!�����rZ�K�J��|���5t���O��d�գ�e��d���?�N'j�����l;�~�B��x����}t��Z���vrj�xz��+�yӊA��>�R[V�/�ʝ��K�M3-�'�����[.�@���e�8=���:TL�Aދ�l�z���AƔ��)��	Ke-��-��i�����%XE�&���BMw�^�-�?�8"E pa�7�Z�WJ#츫���>}^�֬wa(1h칻ӓl�����K���k����V*
gL
��	/�A D7�fc����R��{bt]Ի�D���Wr}̏�d�J0� �[�\�A��pd�ŹXV~��;Q���&���kp�F8��k��;܎-ы@�|�$�Hi����{����1�o�,��( �a��[_(��p���q�f� ��Y�}�%�����9����D� =�%����$�Oڶ(��t�7Obř��,�p�$���i�#��&�s�:�_W6�K���g�Xչ��4W��]���/ϴ�Ӧ��2V��G!�W������)~َ�eG,�000���;Ӄw�V��e?)�,U�W�����8�	��If�.E���,�k9{	Q� ���)����A����ò{%P�Ӝ�q���CP�k;�'�<%&����>x�1/ֹ�͠��@�"���E*�<�""�H��<�2��~��o�����Ư��/l���t������6��d��$~���M�i�= L
��Y������]qDGh���� �ͱ��,��q�2SeŘm8X~dWg~��A#���:�4�lC*\�^�}��I^��1�&����xc���G��(�v�R1yr�x)�M�v/e�O˘(���2�.��Jj����9�|�Z��������~�<��n��S�کz�z"M�R9����u7����I���ټ����|����d�0���{%�o�-��Ds�cq�Gn�K����x�Cթ�r�V�F������q͙e�7r �z�p΢��Y�F��[�o|X��(��u�?5�v+�����6���<��(�wə,�,�%V�Za1��o��<z��-s_�A�}��$g��Yk,���Z�4	�Z_������z�׮��q�K´�Aݾ�{wMJ�)�����(�N����Ki�A83\��(Fvv6򿲦Ht)l@f�74|��a��tv�c���tc�a���Nt���h";�8�D�ы�?܍Δ+��A�K<�2,<<��X��K[�h���4s^�	�K."�Q�?�)�ᥑR��h��1Ѥ:<n�a�NE���B�lB�]J�pE'����V|%�u�'��D(A D\���-y7�R�N'?>l	�=�ߏ����7w8bP�PӺli�0σ#���u�kuuu1��#"P��4$l�y2N�nխ+|9�/&��e!�&������w�b
n	��ѥY��2J�� �;�՛��AՅM�(A�MR�l0���9����P`@�.�k��r�؈�!#��U�6+MX����"�����v�F����NùyWw�}��O���hk�PI�׷�����7���\B߯ά��{W$���&z�~H�[4�\{ܶ6���[��z��8�
R���E��dثs����	\����ӊ+��ݵ8�Ā��F�2���'��	�t�Qegr�,��]�}	]c��Q����(yܢm:��#=���v�1���,<C����[{`��hf�T+��v�[��U�xy�{IΗ8����
���Υ�N��_��xeJgLr��F�t`�	j��v`�n�[���<|A9����|��l�լ�ZC�r�U��R�|�5�p����b·��X�F��A���+z
u�$�A�W�K�'Ӿ����P��u!�-<¦�a��F���͹=x��A�p�.Rjx߳����	�@et-������O4�jV��Ci�Э~�rB;22Ѝ_x��9F+k�<ezC6�献��`ee�����?M.ά?�"H��f�2f�='������e�c�'�����7�]
8����Б�?76.>�Ϣwٍ��[&�l��_1v%�[�4��=�=7MS %P	��<\"��Q������}N�80���J@16S)��{|���#-g�w�������MшI@ �;$���m��-�@�m�5�������u�5~����q��L��D��1aqq�"nPY'냭<�n-���'�h<���\��\�	/ا�|G���Xس�/���=bf��Zo��r<�f�3��l���t�3��TY�p=�@}��/_��7�GJ"��X�}�A��l~`�V��rM|ǽq���J�b=��>I��T_+��xq���P#t���v�NXm���T�p�_w_�BO?K�_0��iq\������)_#���گ?��%�]k�>�g=�}�6^��}Ky�*�I^�Q�e�Kڸ�[Z.�W���"��{�E_UM�G�O�طV��B3F�o�2������L��^��S�
�|�߳�d��k��ć����6	�	 *�^`Z��AC߾��C̞�t����ց� �h��:�Z|K��!�ʗZ���p�����R��!�恊�Y�A��"-�D�V���4!�WT����X׵Š�p73�N�U~+�ȶ���fk��^#(!��m�a]h�:��Y
;�`v�%�R�t��N,.T�3�J�l���k����|Xy k�2*�A�q��;K�5�����٤�(U��4^#A���+AYr��r�ʊ�'|��
��}�����דo�m����m���hjjf���"NoS��iq&誶?2��8�
�Zyy�G_YU�a����B���SK𓱌�*��}�lu�a]}�p�A�E����7	��t�x�F�,��A�߱�4�$b0�ӫ9(�y�����a"�<�Ѳ���Rw>_s�>و(NqG:����� �u0'�t8��1������8D���*Xk��^��?����P��)�K{��Ih�~b1N1�/s�q�9C)���wr/���*So���`��Ǚ�E�p�I�[	�o��\��yK�����'�m������>T�t��tt��$�lǭO&�Oc&�-��%�Q$�` 9Xa�b��f���S-�n4~�9�9qh��������I?�a�s9�_���W1�~U~k�{E�,�󑉾@}N��qKz�aU�U��VH��h��|?_ek���.��#�$�n���%$`�'��4uu����p��V�)P4���ckY2��T~�|�n������߽-<1EHO���~zb�[�?=s+���e���e��oV�H��<�<��Ѕ1V
Ԙ���(F+��VS$��hv�Q'�o�G�O矖����A�(����\3c7�n�vM�<��+>��@ˤ8��������Zeki97H�}�t|�d�ړ2�2�8�b�!㯓������H����r��jx7��=9r8�A%]����+ue��&�K�]`@=u���3��E��R�z�����7��lI�T��퉵t��z"���<�_[�3�T��Z���ꪊL�AQM�PίTCߒ����ܟ���EZ|��y6�z��J{�`�n�	魭b��_O��1vӂ�W4���ߟ��� �!�_v0	*�fڧ��{�Lںj����i�xe��U�E�����H�i�v��\���;ܖ�2�g��n�uG@!�׳>���[�¦�E%o��φ�Y%h!y*�$��]����;���O���$,%%�l���l#)|A' 3�7�&j�4"�M����y�����Q��Ҵ��C��+�ϊ�h�Qځ0��G��Ǐs��v GG1C�wv�u� ��0x7d	9_��	��,���� U(���㓢ʂ�'�Z������)�����qD����&�E�jZ���җ����t뒼���'�x��81Z�f�o��On�=���e�މ�φ.�߹��?���
M	"3��n�f|���=^�=>�F;��V������k��t�������DG�I;��'gQ����d��RRe*vSӓ�V�xq&��X˿xp��e%1û�|�0]��akm��6z5I5���QNG�~�DX.m
�9PpO��v"���Rr��:O�gy?v$�` +�
2����6�4��g�zO��=�4�vD�Z�#�.Q�H_Q	���9|��;6v��� ��(򲞆P�h�W`�vˑ,��^��.��Χ�w���ј��K{����6�����W��� ��!	�ό��U����D�['��Ϟ�/���h��S��|C��f�
�s��A��SJο���Z��	Fs��֨���)���ۗBߠ��4{?�~�X8Pc⾽����᧲x�]��Y� �%MI��fQ�&ob?ֹ��f��{�����M/��a�C�C�%vfE:�\��$:�վ{�Ik���UK@��x5��H6�|�c36��a͵G���{u��v6ub������4Ud�19��]�S������BL>hrۣ�Q���K��{�ξ�!HGc����@��Ǫ_7������iP�y6��,s�h�wC�v�Jk\]J8ޒ�
,n&*�m��������I�j�-�1��C�=�c^��YO�ҽjLqY�	@C[���z'=4IbBƦ�7���ܺU��gV��ӳ�ŏ��L��<�Z������іKƜa/�ÿ����"z��抩UV�5N×v��去�d���q�f+���l��\328���/���k雽G��×}�Q�f٧s�pK��XW��V�N�{�O�+�xkg}�h�mD#��I�P��׎\e�-W������m���d&W�$��V�Ņ�ʂ�1.m�n�)��T]׻���\�@?3O�W����k7l��r�%����_�����|����/dP�����B5Fp�)`�+��U��ϯ��>$O!�7��o*�\Q�pUwF���o2��8�#6��j�HxkC��t�ٌ�F���.�C0œ0 �_\�����1o<��N>���d�FI�N۝l�
��'��r�;0K��-iE��j�nS��:�~�֒�/�A�]���=uU�L�4��r݈�ԴJMJ�R���o���C��e��O��#���Ѿ��=)j�Ўy\n;\uYMj��CZ�1��(�(B$)��/��)0�}s�e��1���Ҫ�O� /� ��?!�y�p�3����+y{k	&n%u�Z���ߒ��V[����O|�ۆ�VQm����X�_��Om&�S�.�D���'P�K�FO� }���Nb����O(�h��{�X�pey|A�jNz00՚�wxil��͟�����#�TK"�#jj���/ӾA��e�z�j.�k۶��(�]F܏l�Ǔ݋�*�A�=�(Ą�# Vo*�kg��-e�� ~r��"S�oD�C�{E,�;��.CP,���Z��X�pw瓤�]���ة�P�H��EJ�h�t��q�g��~� O�XM��d���FV:W BO����[���̓{.���4?SW.12|�_9�v4uA�:��q���J&~VZUw���Q�.�zց-���8g��=�Jy��Z�<~��!�H>�����X1�t
�N_I�h�Ѥ|����⾋@+��r5Vh૰oH���aҫ���Gpق��犯ΜaJK!+_�L�ÿ4X����U�!/q�� ty������Ywh�r���BXfY�O�f�l�����i*�H�@Ś���}�P�:���cςH��⊱\H4V;`m�� �%SV�9�"¾�2n�Q�~ikw7�0���4q �)�#̍z�3KPf���%Şr�@D�u�R*<rtI�t�H���ۭ�����~�f29c���3gT����;�1Mi>�o3r�� 7 �b{G]d����T)[���ߚN9v.}o_���Ћ��,��_%	�%��4Iߖ��^�H����7׏�8�Z�R@<�b���J����Ѿ}�S/�>Ӄ��Dh������`#7r�
�W���@�&Hq�G�h[$��mߟS�W0�ɂɬ���6 S.��ݩ8b�xGGR���쀌�˶����5Ԥ�D�~]��IVX��G��~E��-�m�¿��h����CB!���|��..	n9��(�zGI���_7��֩eE��;��Y�"a	����2K�⃽����t �PO,�As=Dd�|G=g��R�՞��$=.Z���H�@�s����m
��q�����(O� ��v��b��AB}��8l9�;�&��������5F�>�=��3�Eŝ7tNZ���|w��H��W�~������[�3Rp񊉉�!��6I��O����Ok�U6�I^��'�_ܒSyO��������i@�Q훠�
�2��c��n�%�
��:����zj�b�Ne�B�>�?t����?)C=├�ʚ=����wnm	љ������2�)a��D��d�x*�M��X��`xtiIAG���]o�<O�l��	��`r��j۪���Z�g�Csp�7�ϋ$��X��J<�ڂ�J��7��,��i�����y�r�|�촁cF��1]�÷D'T��/3��?��r�|��i�۬E�n�����!D�vԄ9��X�))�+���6�>�]���� J���ς��F��'c��z#W+�KO���Z�C��J?�̃	Q���JoˊO��lj�7��.��-�Ϫ�#�{bPR����G6����]G`��/E�>+VL��s���5{:�uvO��l�Y��7L���aa!Q3ir��������3dŏwhg�|��E�z�S&�%�m�Qk��(��nE���F���|1�������B�4=�a���)ڣӳ����%'
js� �s��<}u�H'C]˭�x�$ǠǙ5Z�q[U�	�� ��f&Gr��> ��:�����&��A�2d�&��n�&�3Գ��ڟ��O���.�s̤��ua]3z���S@��L����<���_zvۑO����y)��&WGb��K+� �ܫ������jX�I(�����Wn�b��_ɩ�������&����'�o_��N�����?"�3�Cy�xAuʴ�:7Q�&�`c�b��ќ�d�E��bl�u~)�Ɲ"Q�`uΧV�7yJ�#0o-����dV.�wjD���2�<:�@����M�֝3[�x�_�[�Y�͑�}K�WM����J�1h�]M\<|�9U���$��DY"��;,�N���S�wo��,h�o�*Y[�A�j�|�LGF-c��~���X�qG��h])'5��� �sEsv�n��"n
��\��ȡ�߅������֭�AWa�û�6��"Oۻ9
�? ɴ�����#�����@�(crq��f ���|e��ݽ�.��C���x�����3�_�J�'��٘cU`y���
���sIM�\7w�9���~�	��l{gzj�8�Qʅ��ޕg��`�G��М�/���B��F6=��N��LbX�FP��;P����8ϢlD�뽃�j�Q��5מ���v��i ޱL�ѮF��v�G�<�eT����`�α��?΂��[=4ሀ�Z����������F��+Y/�������n=��V��~�q��?8�]=̏��+9�6���o�ll|�3�+`�J 6[��ߠ-t��IpijG6����h�����v�>H��F&l(C;8#��R7O���4C�����l���/
'Z�7��㉷w��m�,�1�I���1S^f�e5	���훉M)6E/�Sl����^ :㳈�Y�G�21wH��r
���KIyA��(DDԎ͹�Սs7�^V�o�y�EE�>w��T�~m�0M�ڮ��,I��O��d����G8�I��ƫ���������+�5�<��2B�9��+Bו��(�u������)��\�C~߸t�O�#4<+��r���#:)���M9�-��_��qHL�-f�����MZ"C3���KqȠ�Hе�VS�O��O�ŝw��]�}BbJ�F�&
��P3��M@@����Y�0��!9B�Rrxaa���Ǧ�Xa��X��t���gg�|�ѧ���l��s�e���/��~vɫ�T7y���TH�Є\���cF63>�q�I�|��;
�y�R��{B@��*�����F��Q�<�w�Ґ�H97v�d����"�Pb�l�����S��}�O�H�g�o�^d�����s�=ܘ·Ǳd��e{��3�H�48��B���IGҭoF�`���a������ڧC�ˬ����#OB�w8ޱAV4eВ���P�K���
�Cry��l^�r7E��@D/�m }�[��7�sl��9/xI̓$M���V��i{7�LM&r����8�Ο��Xj���&��~q��~��k�a�)�7@�S�;�k��;MfL�UJ��r��͜�E�z��|�)z�Zڸ�$`�h{ႃU#��o+;i��ޢxR�7_��jq+��hN��'����-�T̟��Ӊ~]u�.�L3��G� .=煄�-v�D���V>�[L<,k#B���~��Lה-��K������@�(�������}z~mwzH�zgTt:y�H�/>Fە'��^5�%mR�-���A��#�L���iK3-�	��=6�q���4�=c�M�YɣFW8��!��f�Ա��G]����^�[�� p-��h_Z������"�?���m.#k7C`l��0�O8j` 7�3l�r����}fv?��Bz�}��j�;c��%/��[�cs�\ 3[�W��͔�YP�?U�C>vڤ㨌_Fr����<��1p��5b�̳>*���wh'����r�x�!��t�h�Ĕ���̇��(��4�̹��%��nV�s���?Y&��k%��ʅ��Y��$�џwѶ�ؕ>�u/�R���ʎ�������}d3���)<��`3��X����X^+F�r���¯.�>(�D�ׯZ�D`\I0��>���]_��?x���R�?3�2��~�U��n&���r���~$ඝG�`�*����KbgX�� ^������IU6iy��"���zJ*lD��oc��� �w�`tm��ӫ�*n����k�h�+�o�lhԬ�ӂ���wA���IZ�P�����%�=���?�t�������k��2Q���a���E]�v`^��H�b�14ai�V4n�!��]��"���Z�]�\��d��J��<��pM:|��/l�����i���뤕�&u�&]M�@��N���ܮ��%����#b��N�6L2�'���C�%��%5��0D���z�u<�������O�G�r��� ˦Hɍ7�7u�j���g�>nL���������8_̇��Ԡn{o+0�Ӝ��n��ӳ=ݻ*�����/�J�%��	NJh�*"��b��y�	��#A~E/禖�ѕ��U^7���{�tG�\d���wv�6�y\D�Y��g����8�
O�Z/7��x�CD"��ҙ��/����?&�g�M�)^�E^;ƞ^\�+�Wi��q5�ȇ������~�&��d���^=�9K�6q���o�������ہ@���Y(B��X[L�"���Q|e��R�����i���H�G�1��N,BX�̤��
8���֤���"� |EA¿>�rF%qiAT5��!2�Js+�� 6/����a�����wQ�����\�|���1�u�6
�\:܅7<��vv���g�Ȱ��@>s�=�4�z���na����X,�Xdd���������ۦ�?�E^L]p^�]�h�F�rU� sn��8���Y#�ٓ��T����͚=,�b�X�!_��
���ӈq�_�x���z݁��xV2Q�dg�m�ۍ1��ņ7��	�K)�w�(�1�,��zGNJ���kz5Y�_Ts��m� AKt����)��[�)��d!���yg%Y����J.�ko���޿B�'���ݒ����}e#��K;���y�ӛ�5nN뇥�itM2�`T�#�꡾���,�fBe�a���񸈵v�����H�8
��s|z�C���(2��i����~TAAm�/�v�"M-�b�
�������.�L�zˍ�d.��:���?�pc2?�}�F��G�>?H{�N�H��$A���h��p�E��I�-��4cP$��Ei��Bz��6�Е�N�W}x��"G���\�r����܎���sKZRJ�B�_AGI	G�7��~���=�^�Hx�Vth2�u���<guNg��&@թ�x��|N7���Hx���=�?����
��AQ�	����W��!��!_��!c�us���Z�
�bњΣ���|y!\*�n��E�\��8/>���$��2�)��%�VL�2����fl��]�XHv��{�SWp-� @Q\n$����-צ�cL27�r#1�3Z왮��aٚ��Ә�R�s3v��o7OV���L����I����M�A��᷶3��F$�2E����_p��x�':ήȄ��x/e|�Fȿ_-mkb�?{�Ά
k��-�T$D&�>�O�~J�����Z�uާ7��pʪ��v�#r���u���l��?�Y��÷�w�.Gs�q6��������m�S4�S#6���Ӻ���K��"�7j���pX ����K,�5ۈ~Gh}�7^�(�b�!����~`�YyJ����JKY_�Q]�Z۶�w��]ow��׷��E*V���7�.c���-B�w]����"��HdS5��7x�"X�!��p�B/���fI�sW�F��	����9RMHY�,�l�����K����/���h"����$�L5j]]����� �	=u�����2-�A����ם x�"�P@.�;���J�q̭�/.ky�y]�]��u7��O�4C1�Ξ-�615���y����C�ڍ���D����=�u
璿����v���=�.tP��Ϙ�SGP;����j������w�c�H��/?����G��{��I��"͠�DJ9V��cL %_}��o�|���0V�Ɉgt6(�okW�#��y��;�Q��H�����zY�Q��,�{��b ���X��\�� ��+�ǽ�U�=Z�1��N��!�ۺ�B
>Q�]$u,u�����Y��͕��6E�=���۱J{�E��?�?�z��"M+���eU5u�4M!{��m7��]n���3��K�,G����4�A]!y�@���nT���z�  Om؎�\f{/�W}�O�}���0�"��x����u����QLVQ\\�]\�y��|��rp�_�:>wmr'[��Jc7��d��O�"Q�����FaZwB>��r_��1u\۰�M�s\N��ں���;F�?e�"0�* $�Cw�3={]3���sJ��mgY2|a�a��-��1�Q�[>�9E�g�d��"[������ͬ�K��b�Vy��S�b�p��K$�j��I�w������o���X=���fp9�ܭ��+K���)�(Q���/�4�!1�ų�S��;T��G�!�������fo'��>B[��Zo�DNl�Y�!]w��78��<D������5~4!]�4V�
�CH���$�DM�9:Qq�Ȋ��T���2x��Ĕ��*�:7D����c�e�Ag�f�f����-RNd����]�M��k�&��RPP�EW����"J_��x�X������}�ր�\F��Y��x�`�L��1b��l����sB֋&l�!���qTi�bsn��E-]ُb�転��\�O�->LO�n�� �
���{?[��P��ߞ�?/I��2�J:�K���۞ ��)��$����JT�ݯ�p��߿�V/TVV��V����h_
l�Sa��e����aX�#C���T|޲�@�ė����R�9�.��3r�R%�b�@�������pϓ=��f��7Ѽ�5��H�!�L�so����c��}0-z5�Ø	@��ӭ�+Y9~���ֿ�#��ɑ/�.�Ӥ�;D`�QVьWei�q����°�&@
t��D;��4��S��루[�=c�Nο���6]]=/mb+���V���)�v8�%ϫ4��F�:3�[��ʬؕ�M�9���%���jQ5R��g�F�9�i2۝��9�H�c/���lJ�o�qA�pX��kl��X����5���*�_(VM���}g{�L"fo��h?3U(����.�\ɕ��ęA&��UW�0ZڏO�0o����E�7�O���p�:[������x�y���'9G�2T�K%����N�hǀ�I����\���@A��~���h�P�=06���΂&�]]�ík�1���h�;˧��^���5t�b�[P�l���lt�uy��a+�R!���	����F�Ce��S���~���}�Ac�`�Q��4(U!x~^�yrJ�N�*a!��[x���Rxz.�}-��˵/�D�ё�u�Y�Q���bP�0����-��G8�'rZ��G�o0�%=� �b�*K8.$j�B.be��7�5K�7�t�[��j� ���"PX��&G�xvyޣ�%��q����ȁR��VB�	 }�B�E�M�I�2}�����)�����Yj�&n"@�
��/�OQ��G���v�Ȅ���9�H��Ô���X����� �":ڛNDM�Nܩ�����B�+��Or�>�u5�^���콝����m}�\�)�z�
j�==��p?��ю9�M�ixfϼ���[�~D;��I�r���'�-^i|ړ�������ܹ�J9�'���u����r�e��ގ���S\`Δ��P=��W
u�$-��纹�9*7{�c�����NNҷK���t�q��t"R�m9h��Xo���_�yWbsg;�DGC#��v�L�t�>�H����i$�
݀���!�Ə�c�:�
̅�,�������`�Q3�e�9�.������+)���zVb�i�WPds��a�� kyO/�����W��?lX���a�7]�!cԔ����//%��H���~���r7Zۈ��S�axA;�Y?��o��޸�-]���j��ݙ��4r��SQ�����Ȋ���@�ٗ����C����[��F��{Zܜ�x
�0�rL�}��Dv�jnn�(�� V^p���j���\�W��.�k�팤l7��:����8��V��7��BҼ��:z!���dO�7-_���~���-�9p��AS�'������x&5a�%+/�?��	����86Y�H���,c��y&�c��U������?�Z=�u�)����}3t��;L�^�Mj�xk�L�znZ�R��wF��HP�h��H�,	a)Y�?N��V�xљ�[d�絧��q��B�Cdj���J�4ި2�d_��igU���P�H��� �t~�.m�5uZ\6��e	�"T6�~��r�N�έ_��@޳�R��>cmmu
�u�=(��zbڑ���<}t߅����V��D�7L�`r����b�c��".�ZX�C��~� ��~F������H\��Eʌ��T@˘9�=eA�y����p�xơ]_wV�x���G=+��;�u�nɨ��3��U�2'�E�	 �E;��)�|U�5fU�#��K�0:�jj��%|���L�E;w�A��P&)>��w�l�iX�d�$R���>/݊ K�q�RE)#C�W�\\<�|��yx��>ѓ��V��f�f�X�5�u��5nBBͯ'"�k��1Dl*����;�����ι���ݝ����ް�)�5�@��7����\�|ȷy\�&����i�9�����ʎ�Аp��"�1[��H��J��E���h!۹���pq3?��~�|qz����t��1�Z�D�Sj2�x�꧀�	3���h������TZ�α!��7��矿��1I9\����u��<��x�����>C"grL���N�&Y���-b?��ES�՘"( :�s{h�B�^{�3�b�"����iNőý����C�K�PaW���_Q�?��F�� � R� H3蹹��0��[IUCLK�zb�:���s� H�n�^f���2���+��:�j 1�Ƙ�B,J�'P���_?���O6 8���������k%b�X�~Xv�	�Ri���--lR��E����[91M�l�GƟ1��X����\�����Wg�utB���"Z|)61ָ$��L,�ʐ�ay���f�mV������Re�b,Rbs����$˭���$���&��_w��qq���&��Xj��@O����l��8�s��$���8@^V�L���{������%�#�1A��y�OɦL�7H���7q�o,Y�~fe���>�+�(m8����qZ̕U��Ц1�d:�L�+���� ���~h�^+�$��D�^���h^�t�9��6��;��q'���a���vUc�6���Ѥ���Lz�:"�2�m��љ �}���ut��M�N�����]��Y$]\?���gp�)�S��X��ωg,�%��fŮ��Z��V�<޲�BBBJ��C�[�k��]��������ՅkgIԋ�~�ʆGΆ�*h}���&��M������( ���k7CNóy� ������yu���[�ɟ�JV��8�=u ���@J�'No�b[�o��j�s�#�D�V��j�&�Tq.1��ºw6#N>���mA q�o�^�N��rOw�r�"�;'PJ[9�K�.�{8��>�m&��z�Z|D4���� �O����W#邃 ~(?���>�&g�
	;wj,�~�:U� b�<I�A8�SW�~�gd����;4���Ш�Y`��H���/g�}�e�Z��p�O1��ߒ��ja_sZ9`XQȬ��84��������!*TunѬ�����-�lt�c�~�E���M|�ؿ��t���y�����Z�X��7� /4:��2�[OWu��Rl|)G�Q�8(��A�s"�/:_���K��~U�����=r~]������?q�ZTpJo�`�)}�{a=Ӌ�P���s���0L܎%�F:���C��$e��`aSO��j�è��X��ߍ�i�(O�^<�)��	��y��ڑ����m���G�`NX���1n=2��º�;e�$��N����������c'��Ŀ:fc������:<��d�E[X�/�0�`n���!;��9���$�����"��M�4���N�4�WS�o��
��(�r�)�R�	�f�Y;̏k��^)���^�.�'�#<�)#��}��B
�l1�yp�V�=�C�z�ǅz)j��?p��r�)��a�7�ȹ"����8ä�I��=�z6�hfHX�8�� _�.q����xdn����
I�K�wc{h��׈g�)l~ֵVe���t�9������z��N2̀�9?��/�g����=�
d��QX��z'�R����][�$��X�=��k��U,�~"��
�5�N;ڲm�ӝ.D�PQ�Gݠ���a�+���n��ۃz����!!�t�)�:��^��3
���kϒ�ω"(�zC.-��PU�g��*Wo�n��O�ut:A�'2�(�<�=������swd���'�ST�^�GJ��4������� ��ϬJk1�1Z)�*�g�kOZ^�B�����Ѱ䃘y���"��8�y�<�����؅��d�Z�4�/�كi2u���J;�C�ª�U
������[��W\�u�~���V(�w���AOA�i��������f�
Z����\U�*l��};C�U�sVYyĔ��u�;ӽ� #���+��Qz��^�J ٶU�o,�}C`�����A1c-T>��L Ɵ�������_m�=􁌻���T�5(G�*]�X�?�)�d���a�M9�c�z�x��j��޽�ȔaBݷ�A��o���F���K���0�<��u	O��ĉ���k�fc!j�]8�#k?��y�&g�m�O�%�2^cp��������ŋ4�9����6"��ӭ����Qv5<��n1�4�s:�au}}��]o׶Dtpwwn�]C��]����N	��������[p�`��{�W�U5SC�ݻ{�Zݽ�y@X����D��!ޚ��d#{kK���Td�ol;�d� �����#O�/W�h�k�����(���{MV����m9R����})O��SΑ/�7uV> �������EB���00�?u���ʆ	��p��P�ud,�P�l��~mq<�`��[7���HY`�0I���NQ`h��(({�Ȏ#~�ō�c�ۨ��󻇟&��zh���s�Y�`�}��;q�������#��=a��F�e���o�θ�e34}�4?�\0�����O�9�́��Q�������J��iY���\����_�Y�A��}��6=��op
��2�1���Y"e���Ss���i]lǝ=�l)�f\��7�i�_s�wUNC��dS�蔚ܿ�'#�YE*��YUnͼ;WgJ�JU��~t&¡u�[��!q�2ȫ���9�9~�_�-���z��`j9����PA��|��+V$N�rJD���A|�d�y�>O3L�+Û��Y}��q�g�M�[�k�5�o�r?ܒ5�O�Py;��R�[[/����(����f\�����َ3,��r\��m����� �Qo����?���9I�S����{�
��<� tG����]S
��R`y��7�K`QeM��"��?SDn:�J��}��>Gʌb�=�b�H��sΓ.���W
\�1	�_���Ɇ������=LF�����Vʚ������X3�%$%{��B�1�C�m���*���XO��d<^�w7KR%nvC��(�7F������.���ô@���>�J@�$$�|>�0c���H�&��3��4�$/<�A��"�(�&cը/���]eƅ���=���Σ� ��m�;���W]��������[� e_�{�]l'�u��Mgn�s���wJ.���w��nV}��w�=�Q�<(T׶;��9W�.�7���}
[�TI���U��u�R��s�����噫�t#w4	s~,�7}�� �?P��%o]���3/bWQ�}�Dqu&��U����$y�U��st�����U��/��J�6�=�/��0����\t�ȓ�v����ˉi�Q�շ�ɢ��}�[&>o��DV9�w�O�+���H���zS��\e�ݺ3B9����'�|Y��D�2 t�� ��-��#G��W�.P,�;�1�;`
�?�A�u%�'������+��M�}�c�}��J
H��������-�
n��]3]H�����s;�- "�����S��'��YMU�e5EUx�}�"٘�(�\qG|i�E�čv#Ӣ�" �u=߂	I>ɀ�ԧ�ާQ�Mÿ#��v�����!X�%��+�8�}������&��n��$�����ӓ��2-�mY��㨤(��RbvŬ�(����7O�[�����#H��z� ��9"�����3z��O��Ipol�����Ɠw;�vNf�曆�;	��Q��W�2~"M&@�Ǹh��f�&Q���-���{�b����¢�n��8�@,�s�r$�޾w��^vz�pals�r*�C�Sw�� ���U�Xɓ����z{��zZR����y�K�����|� U�������Cl:�5�32�f_#�w�`�$���}at߈w\�o���0&����̠l[Xn��f�> �B���QrA�P�c���bn ć~L3�~�#��7�鱕�`ii�8��9{�x��]��Q�Oߴk?�L˟ J��1YA5�Ү�+�+l+��)_��cG��0�*���jD���bO	�"�Q��7٭/�rG���JM�ir4=�C���4y�$�:+8ߞI����?˞a�ahq"5/�}-Qfs�^��*�l��؉^V�2�a������9��Nh]y����<=�o�����#H2�Xr}ge���;������&k�w�O�'e%�\P`P 2��ab�Қ��/w[��r�^�;�[�l���;��U��Q�;�Q(\�E�U}ϙ4��p�Ȏ�O����5����&#�.��,���Y;H���C�F|�0������e�0s�B�f��9�Vw(��`�1��'�A�n�S�Q��b�Av�m;�l��oh'�v��yЋ�9f����C��9	��b&j�!b��cq:��A��pr��� �ja�+W��/8^����_l�D`��yD:����M2ұ]E��ЎU��뛼�F��X�U�(ɿ�x��g���*�@�ͽ�����M-ͦi��
=��7�ꔹ^�I*[�K�,��k�X�����?̚��2������Fo>*--�DF���bp��i�LW�LW_Y����ߛ��Iג@��na�l�+V��jo���=:����`�(�)�Y&�=�ȿG]:�H͵�0�f��#����'.�c'V��K��! ZtL�'+䄃�t"Ҋ�N
��l?N�eD��
�c�&Ƣ�M���+>8sv[g�t4�}4Ӈ�j�&�ǵ�K07�WT��>��5�Ǡ��U���D�	��"W�c��y�� ��;^4p��v�ù9�7Fa/G���
�3ѧH�C�0��\������ɋ��{�n�輳�`s��%�������O�M'
�{"ߤN�d�bkr����&S^)�����q}�Aql�[�ȍ��^0Qڄg�?�i�O�����Р��%Ǫ9�k|ߚs\��!8�M,t�?c7!�~ۦ�zr�d�KI�R��We�w���4���^?i��H
9i�2�"�\���W��_�P�G���*<�_:��- ��$I�=�7b��M��*�}D��:l4x�{�K�%6��xh5r|'���2�g��7E�'H	k��b�5m�y�VMj)ws�0�� ��l�~d�âj�8��{"1��H�-�FaHD��_���᎖g�˩x�K_z���Nn9d�d־�lPr]�����3�0�!�Myܜ����`,�,{�f*#A���/%� �}��e�)�D� �H�}BuSR�����Y4Z�uOHo����6b��?�(gÐ^���_�j0���v�"e4ފs�Ys�ͪ�-g�����{CYI]�bc��2i��w�e�ǟ���!��F�������7š��۶�߀E
�#2����ߣ%����O!&'3�#}+ �UA�MMuHH4�ú��풳e��
�X�'.m:���4p�̻IBq	�����'� �$�UZH���VK��o'Vx>]7ڷ�~_�L�s�UY��x�N\x����+qY�
���{���5����xӼ9���]y��ѿ�X����L�m�+�o8J{�	Q �$���YA��|x������z`7��$s0�6�[�=ì̀Aa�Mt�R�x�*�!�;Î����L��"�Id���N��!G�ֆA�`G��Dc�������SGF3�U=(���b�6kMwV�M_���{ ���9,��j4̚a��E"��B� ��0��L_�N�S1���*=8D?�ӑ�}��x��|~._\�-Hٖ�m��+ω.�I_�UOf��ݙ-T��P*ѾD��&�{g������RF��Ѕ���ˉ��?�.��p8&�E9����<�!4�}l�7߬p֧^'R��"�5|B0H��9
�/�Il�6(!XZ�Y*d潱V&N�@���`G̱e)�ʌ��R>hLf-:������l`[c%��ĥ�5���Nk)d��J���#b�?R�q���&x	�fxrJ~k0gq���xw��q�TL�ψ�Z� ]�t��gV/a(@b|Ӆ6�$�dm��m�x�#��h�4)·�ɣ��N>��)��,�=��- ���g!P��x+%n�V<��qPv����e{���^���CkØ�f����0�t�$/IfF��'�ҝ@���g��	�ˌc΢��`�|���7���ǲ`���J��+��m�n0���O�9�@��H9)E!u������_��6ÂȬgIO�n�үΧg��m.X��Zl�bO|�Lfh�(Ͱ(�����JK���V`l>�W����j��G��w��7]��mV�q�N���Y;�4�Ղ�p�=���)�������?N�cbd��1�WZ�O4�N�������k���b������]����n��8_3+�mabp8��\�OY��@���o�T���蟞WR�nj��|!*~�yT,������ζvANv��jC.�yYz�D�,�����:~�6k`R0A��u�-�K
PNB$%.2��>�!nP��Ӵ���wB�h�<+���mZ9�@{�<��Ds����Z�6z����}�X��u��:������PI����|M�?ʹX�J�iI�"��ſO��r�w�9�K����ws'�O��$�ڭ�D9n�n3�%�V|��V\4�mO������kJ@b�J�e_
<����X�����F��P�
0,6~�D�l��� r�L��sYAU%�� �}�h�	!g�ɦi?QD��Μ{W�#��2
e�9�|5x������9��j�V����s�j;Y4�֊f���'!� j���G���b%e�5D8�u�UOPUԊ �����I��F�wz��ЉCv[Y#��
�$���6�k����㶷2�����ovB�-�o 	[*�߶N��/�uEOy�u��禑V�u7�v�˟�9fy�S~����"I�>� �7��P;��>c�w8����K�	p�]�̸S���6�����ȣ����䜃�2V��f��ࡏ"!j��R�V9���t���[א�p��V���^n|~�LZZH� ��Ǭ8-������zU29[$a[ET!,�G8����ec���r�M��DP.�"0��7Q���"�Y$��H/"b���N@X�-�J�w����Xv�Ǐ�(�L�����u:>R���$�k%p�T�}�����s_�]|��q�l����qr4�������s��%�r���D��猾V"��nʘ.Qk߯��ܹCʤ�;����p���Ws���h�ى�YSx��[�l�?��Ln���rڮj���sB�F���3���_�Go#�y�6�%FcH�9���m�
E@�O��1N��k��C������2��X,��ܮ������7��ſM��y,5{!���.%k��a�W��	�7��@��`t�U�z��z�¿U^���k�2�v���6��#�~� �k��b#y�yRr�� �?Y�gOs�m�T~**q��{�i���-����\�	6�Tܵħ�}4@�����z�db�g�����t�����jI� +0���wtu�D}5n��Ql����G�5�y�M<��!�����ڱH7�����i�����?�~�j'�2���V\f����� �T%s^ne�)���U���	�U׷���	�8Ĳ���3���`�"�h���vāΝ%��%�2�7�6D�hc�z3]
�:$����1��:�s&�~�O��~���i�[/A�}��Hs#8�n݊��q��[��D>>�5)#��MR��q�Lשmj2��X�5x5&��F����,��L��҇�R�$�V�V[v�e���N	i�+.�>~�x�ѐ]ѽr����� ��Ұ����l'�Vo��k��Z+��(�]�U� xL���Pf�Ra��W��ͧ|\>��=f�EWJe ��Te�M`�z���+����|�W7����p�F�l�^E�Q~9J��s�V5��}�C#���a��;{o p�{o��a�a,gl|j�#�Ù8��R ˦��)������u�c�7ݕ-	��+�e�)~�ÉOe��
�55�>hU��e��9�;E�VYy�A\ϞX���W8O�nOAZ�ߣ�%�����ľ�iG���p9��B�'ٵ���Hz����O�gi0�1�=�r>�W/�b�q�C��_k�$8�9$��2�; @Տ�A�����x13�u�>�c�&��UG2�����$ݫcs��<!���5<����h�MK �2�~�h͔"%��H���0����ƒ��B)��88�IL�A��$EE�s���2��.�=+D�.�߳������uI4��j[|�>�Qt�}���'ܮ��KG���W[;X����V#� bh=̭S$^l|�c�|Ug|�?]����	DǱ��U�D-�*3F}�?���Q8�aYQ���n]��Л�d%T>��z;t|Vj����\�nф������j�$Xʛ"�ġ����,;݄�o���5:gto���&t����TBu4�l�Dn#[L�EނP�
�Kh�a@���_���"�<�!ZZZ22�~���#"�	�Y%T�^����F��]^�/�t�>��'��0Y׀H������P�T�Xآ8�ȏ����"�/�?��6�����gQ�@�@�3�88�sr��{o\��@L�ZO�d���W��T��I<��1|�Ε��5����a��#(���ܲ�vo�8��3O�)2�r�i=�7v�d�Ɣ����cƮ��ٜ�JC���� �����N���>�mv"�'�lE���j	���#�vn�0��u�Q��x�:�mW,�"�Z��Ыm�ViKoֺ�����.r�1""nC�G�F�0�f78WKX�d�W}%�(*^Y=/��u�.)����\m��@.AM7�Tn%VLJ�_��ɤ̖W�1Z� �c���rja���'e��ffwUו@5$i�T�~�M�>ܬ�u�]����Щq��̌ƞN�J��W�Ŋ�T�RZ�ڐQ)�;^�~��8Ckh�"ĨZ��l
BB����7��3h�|7��8��)��k��7�����R�z|2j80�&����
���J�0bP��.Z��	�-��z�o��0��	���c�p����J,�%Z>���-�b�9�S`6��D��#鉤_?$�����e��R����w��6�a<}���d�b�1{�wk�$CT�����Q�����s�oY�p�N�n�~i��7#{�<�/�ca��L���k�g8�a�!U_��T�ސ���ЉW[Tc ����bP��䄭���
��0U� -u�.�Uk�u����R�S}>�p�&a�FW�>+�cp�GO��qS"i!����L4��M�G#>��N�X�`/�NE�/����*!K`l�Fu� �r-�\����|�ϧst�kD����������}�>]����I���BkЄM}!L���>/-u!���o�fUŠi�����l!����
6�����c�L��ȶ��yUI0�S�5�(�@�	b~}��+%���D>��+��2[�Xvr<��xC�����&�
������_��6~���x5��v��qc�n�p��N[�8H�%��"Qԭ*r�(a�j����z�CX�`N�7�lt��_��2u��ÂΣU�� S��]KB����괆f�߻L�Si��ᄩcV�y-H�3���ɦp��a$$��MGN��{�$0��oFƧ�bz��]?���9� ���@�[NɋV�m�����|O8m�:7&�@���I��(�l�Di){q���_E;)b�H<��O�Ej_�Ʃ&_�Mx��n[����е��s4Z�>z2-N�F�P	��Ǿ�#�[�N�5��t�/*�9q]!Z�<}�~������T��|h��k���T�!�??�pm�R�
�\b�I���!R��`
�d��!R��w�8 !����3�[���ZR�3KnLU_G�B�4�;�l̳��=1F)�c'�_��g��Y� ��Hk���6�H�S���H��r�%� q���aQ������g�v�w-��bN��w�,�7e2ِ˔Q��ľ�.)�B_�����pI�;�����ɡ`C�SR�σu���L�b1L V��4L�2v<�������jv�AWh�F{�wGf�_�Db'�Q`1ZM�O�?�����&�1+��,��X�;Y��e��?�"$�RY��i!�6��Fm� .�l��4E7�xAy�����2��$tt���kL��}��֞����3{�TCOv�3��cS/���k7���'��G<�+�Nꇅ�;,����S_��%,I
���~R�_}��UԻ'�WDϔ��v/��T�H�k��ZTv�D�h��dZ̑���/��t.k�,����Z ��j��#�pn���v����y~��<�-�+�J@Rw��a���N}��a���:HKS�,�#��[x	$Ҿ�	ϸy "���w��wJ�
�c�#�3R|�]��Jj	��|�����º\����TR��ݝB1� A=��-�!�w��W���R=��\3�=x
P_w.q�X�����tvi�ſ1$��wF5LVsdੱ/�~ºt����̜m{N<�K�IXFv���R����lܫ傖W�2f�H,���v$W.���ͨ�%�|�W'2J�x���[��Cyo���mYNf���يP��V1|B�Qn�{�� �ˇ.1o[Xv�La!�Nlp���y���Y·YG��; �X�Ӯ��__>+�Ὅ�N$l�L��(��N���室�񪍚�����kb�B����vlI�4j>�Sp�5�A=DʭD��ƛY�����ϒ�V��Z���Foy�xA2�
�雞Q�0�N}�z�ش4��)h�����+;҅J.$b����Ũ�U���撃����z��s��3~�����{
2��Z�G��>EN�?�ݟ�Y���'m�Wދ<��a U���'AA������[s=9�F�wLQ����MP�M�񻪀�T8������Μ&��`���k٭m|O��:�"I���7JXA��k��&��#�&ex�2��l�/3g$�drU.�f���P��������~�!ɮ`�j�~����ƙ����4�O�e:,�{�,2��_//G�52��F���7r��R6 �z%��}�1�v�;,ڰ�q�sS^WTc��R���-s&��G�&�Lɻ+3�5���r����Φ��7�P力ι%ޠ��	"S�O�A�q�ۑ<��U������ ,%#!�c�|E�.KM[>�m��f�*yvv-�A#�.;�	G�"*j13��GI���ɵ9�
`�R��P,�5=<�z���)s���o}�h�����o�êFB'N�=K�T&r�R��p�Jr��>��[�D��>,���ƣ�/գP&��c^k�	��C�ߑ��\�q��С���Q��-��h��Qo-�yY��
EW�ȱ���T^�alF�}��C1O��rM��u�8�:�z#�a.+H����
�y��(.��V���?��I��H���G/I�xB���caI��0[����t��N�WWϽ��͘FL4���Ť�3c��Q�z Qn}{]Y��˓����8Q��(g�.H�9�rSfXҝ݀���>�۪�\d<|ըn�I�����p���Wt���vM1�@������%������+���	*��I�Q�(8>(Gr)~����W�;	IpR��5�����BRUS�`!���?�|�.�#f��cn{.�y>8u����Z�` �ts���6^@)�U]�V`iI%�ʐ_S������uC���-�v�ߞ'YMW j-ty�~@�׮VIW �o�ټ�� �,gb�鞠�s[��(9W���^�d�$�ǩ#c��_f��uB��0�I�1h ��4~|�j^16��H>�ʋ��J"�<!�t�5�쨧?L� �G�k�z�Uw��ҩ���*D�����I[��$-��(�������֏R`˽���1VV�ފ��7f��\��[�s�[��X #�B}5��`��{9y���EW� _:G�w�%���T�2I[K����b�
{8��yv�ǒ�8|z�9����x[7��yO���(�r%q�u��=B*����g��H����X�5�UE��g2�OI���&0%��^��Z[z�D��+X��U��G�$�����^5��:��KS:J2���̥D�M�+��q<|�I�d�Cl�a�����{�_��k�r�oPd��B�T��3Y��Hn�2ޑT�~��M���,��XV�}�ֶ�!�l4��b��4��R� ��]�;ߐ���>YJh�/����˔4#n����G���x��E��0�얟Qã[�����Rx����<���	w���6��e��Q���G���º�apX\� myy�C��њ��h���������y9��Xh&��:]�!�`�Vͮ;M��C�W�ؔ��s{[>���'z`��U���U^+��n��4"x���X�*���~�.�xP��y��M~�[��2�J��Wm�2�/J�k�OW�	r�"W�P\�^���x�(�&3K�8}
6��:��Y���Q�|~' ��=7��
�\?�������>���ٍ����X��[,��P+�a��O�݉ȡ�C�W#3�8c�w<ͦ�.їV�r���[��1�;�S�������%�ߦ�wbk�~�X�ω6EEh��3{�d�O�	�e+ui�D�G
���� v>]7��[NI�ک}=���^4>*!�����p�rv�L���[G򤢟(�%���d��|ص���mh|+@C6CG�Vש����������_��߶2%T�ld@����tg��*ÿL^��[�o�.�UtG�����Ȗ�,�;�FɈ8=�C�Ay-�����Nz���B`��~� {�Z	������M��T��%�>������g���R�V��Ɔ����P�p���SѨ��hH�@q�ᩃ�E����8�o͔��FٻZe��m\�#��;�b/z%�]ުq��xu��o��o�;��ؒ0M+=�M?b��&+8��ֲ�S����W� �%(˪�������<O��Þ*$㭝���ď͔M#q�,mR�Я�Z!KR�R�gȠC1��r]��ya�&Î*k��1�lӹY�WY���)
��K!'
[s@�6��Yo�+;l�)(��G�1��;h�T�0�j�C���_k��~?+2�@ �$a< ,�������s�����J,�r&[��f���Ñ���J��+��#��zF��~~"B,�O�:��SV	�"7��xv���.�i��?�q-�������\G����,���g� �on�of]� \j��Z0�{���N'�����w����w�.��PPΑ����^Rd��q�P�M��H�)Ms�%L��ڪ��噵k.w����~f�WVWT�7��χ�O���aI��B�4��%ޘ@]�-��|��]v�ں53��DJ
B�燵[�ԡ��!+%�6�'�����XT���5��[�ҙ�Z:׬t"x�5��R���JϳkG���X}ɻ�	���H&���N�n�Ʊ����A����ٍ˩��}Zn?��w�7��`4�i��4G����|��q�B㟧5�滅��&;�j�֘�\[���Z���P�t�L���s#�OI��s�^(+�VA\R�q)fY��vZ��>�y����Z���'��n��I�y�zW�5?]{	Tu�C�����M=��=�k�H�0�R�+~˱����nb�X���JE�CzrJ�s5�7�eaa�m�ǲOl����T"���B��{J�&³<x��O�Ft���ƭ�ϳX�S�U����"q�6(�zhfZ_�lR��z'ab���~��s6������.E#�9a�S�����W�>kj0�1T�Nep�t���B�����C�&B�̖�$�~��gs���!|��$n���ihm� 1�)jg����&�/��#�l�����L���B>f�x^ӛ��� �k
�i��>3��w�:��?[@�^�؇<||�0c
НR�|d:���X�Dڷ���	-�p�t���&~99y	g�jϏ�ZZ�K�b>�/��^�RosO��gB5.�ם�wwkJ�8� g$w��~��j.��Lx�>�͒��hl�����S�W;�vz�C§հ�?J�D�!KI�L�0&�`[-�:/�9��1�������V+�R�vT����u��3bN;���&��iE��WQ[�X�§6[ 3��a�8�nc��,�!	���:���?z7�*d.��}�=Y&�7B����i�d�3"d�AZ��#'��S�/^��]3gL��	����-8I/Ư W�}�h��G�+��]��}��m�>�sr㏀���>D <66�Mg;���é`�FtP	��N��"�{F���bRu�+�3�q��l6�oY�� �L�p�y�,'��MJ|��]u�m�����|����کF+�񋈩p<�]{uMO2�ǁU�0E��l&Wl��&��%i�!k��e��������|�S�]>6M�v�YK)	�n�ڌ�wmmP�X��i���g������pլ���[�'�JZw��.�˸M\jVE��r�΍�^�t���EÂN��pn�ح���9�.h
�Ni2�F!O�������8��f��@id�wHI�V$�Ңg�C���[;�rHUhL`��Z��mÉ��ur^�K Z>=?�	Z�z�<���`&�I�~�E��X*3��O�/U�����r%*�?1��+�7	�O{�_��i��1������}d�U"�5_:ε�vωvQAd*�G�%�<vF7��ؐœ��yA{���c���e���
��k'fe>]3����1!sg�����#lF�
%.��b����N�����?�("�΋�gT?���v�7H=v�#緉J��Z<��[����v�H��hd��RĕKh�՟�u5�J����3����Α�2�@�{w$��fN���8�B�8n"T�e�����zo�⪊�X�C+�����а�EDr%	*��Lލ�t	
**x�I����i���,V�^ɣ����A'm�8�lr �PIjUdJ;�����tt.GM�/P�j�����lH�Ҝ���%�yv�����7�i�5��'��?׎�X�i2��Ll�F=��6�@����Yg�C<��$�p��b���*�yY��'�k�?D�E��s	��y|�rjt2X+��S%�z>R�1Po�sB���k%O(ì���C�P���v(�u��*�w�r��
YcY��2"
2LF� T�1�\�5D�k��0\n���d���I�����u�8��Q��Ɠ�PPv�8�	G끝��h�s��:�vF�S��{UJx��tg������dP_��Io&����o:���������H���r�M��n��-����۵#s�0��M���L&kw���q�Z4L_aX�e����!�e���D�0�<�#g�#u�!��|����Ň����6n[�+r�~�(>Cl�a��a`p�T�|�Fx1fq�	o[�Ĥ��ͱ����Uk��G�{vhr{}k�S�;�ap�?����ڶ:������VG�
���>��"Z��t#@��ز�':Zy�s�U��'��L���ȣ��R}/�G_V�P�F�e��VR$���V%f`wU��z��=�ЅD�������~����~c,̂W�R�����)�D��>2u����O�92�`�{J�#�"��1��\G�>�oP���I�1C��%0���7�)��QE2[����{��~�z�Ƀ	����g�wT�G-��rr�ޖ:���)=�z��5$k�,��GKo«W)�%u|mC{������ 
???`����e�����[�Z�C����;���Mr�3��R�ݸ67�-��ї(��W�j���R&֍��/H�6$��8X��y����"�Rշ����k��gk��6$A�uKk�X���-����Lw�u���Z�2�m�}���$����]T}DЉP�8����_�8o��_�m/�����kŭe�U��̺�D��M&�x:=��Et���_o��� W�fU���*�_��H:lľ����o��`�|�R�\�O��`SCVe�
��[W�O�\ф�cK&8��<},����a��ֆ9�)���t��;,U�n:�Ԓ�C=v*,�1A��+�q��O�nM�~C���:O!�m-�PcH%C[�m�rh5�q�Ow�u�S�N��#l��S�����pYq���.5�$v���6S�����'.�s����O��.�	�����y!��O�?nv"��<�k�H�I��8�+������=B���s��c��:,�~C�^��lo��	bw�$�n���IzA3�o�2	^'7�~��E�F�G]c.��A�rB��ܛ_���/W$���|��^s�k[}���\_zk^9�1,>��jߩZ��S�d�0��8`z��S__?����*�?��E�N8����+���K�Q&��m��nO��`/�eFd�įi���nk�s��!���כ7ĨW�[+����M���K;^X��+A�����]�MV�����/�f#
Mͺ�gR�^��!�fT!�s��q�?-�3�S7i���M���� ���,U�ΩP�"qib����c�J��_���`gGL�(���u�j񸾾�\�}Fm_���� {�0��pd��်�B�VSՈ��I�3�:i�������<~���}b-~��ݴA�@���l GMWnU�=��û���,����pn����Z��O�#>�p0[p�7��1��b����Pf�԰N�q�鴤�#��f�W�\"��y��Ȼ�3�)4r���"�P`y�R�ٜ�3�(�w�w���D���A]�k�X^�-�~��(N���H�����I-+Fg�(��
)���_�;�!/h�%�N��&=�9Y:�k�?�.t_�CQd�C�m�H\�G��`�+�Z�pw�m#�����V�c����y����hȡ'�#�[Wv��`�G��Ko�$u�CJ��KV��S���O���~.��fr���MOi��Y��{��H�	�Q&M�����B�pL�R8lox�Mq�%�L�/�����"���m��?�o<��2d�Gͅ��\@(h�ޓ��1\����$ �m��+Z���ͧ�OX@�;�rmZ�R�&���V��m:=��~!��Dm���L�?X�k~������Bu�]�;��;&��C�2���F���11%	��ȡ{�)��h�/4�W�\bw�����Z�6�:��Bn�đV�� ���N��
�Û�Zy�9sI��	��5�hz~������\�N�g1��k�T�қ�x%x��9���U��kv����W�������q�p�:#�<Ƽ~}��fs��4���P��ͭ_���n��� {��+F�B1\��f��="�˸��x�h�9�\&dJ�/�6� �K�����7�*�L��/rB�$E�&��	��N�[�i�{�m�k�G̗���2٠�72��m���z>�fx�7�n9��W��k4tI/�Yha�z����Ybdff�������E���A�2����cV� ��<�_�K~6���/Y�V�V|��,����n�m���n=�����"{��#]l��qI��)`�ܘ]��Z�7�Qstv�ђ��Vن�+,���(�D����M�2�k����^���
�������A�3���e��WpMG�)�,�U_?�ܨ 8�*o�_�=�B_���Gw����v����s��&���sX�I����є�}~�P��l��m+��'�|�^	��==����ཀྵd/��<׸q�m_%�����zV_O��٪nU�mƸ'�۩n6W�;Ds=f��79q+�ݣ;x���K�f��-�Pس���A,����Z���e�\ O�nb�
�fNr�}W�� s���2���������P,�
��%TX&�ЈvQ�J�gX�'"��ǍRm�:�E���;˶���d�֫t/k���<�������$@��|]S�����E�
�����Ro��Ƥ]�w���%9i�r�~_b-��!�q�5�)�b
�D.��Ñ�ԁ���q���B�ҜCuKfM���2z�ť�!�
���>�z�|\�IV��Y�mB����8�Uq�-?��Qϔ��}Ȧ6�@'��!;��J�C��Mn�;pvwr)�ܾ�uWWc,�3LTY���G	d����%ť/#w�PYSm��h}ca�E����C9$d=ga����[҆�[��2�,g�ce�E^�|]��7Ox�)R��7��/|��M�DS~ڶL�7O�#$"|�>����a��Ų=]���~FcGiim�W��V=���@V��v Q���;�8+�4�Q�ޠ��t�hfR���G�`��X��@���*F�2���|NP�$�f�;f H!���Vh����H����{
���uQ��o��)'�-\��_��X��+�(��E�Iפ)��ɕ �?TO�\�NI[�[Q�ϡ�`�N,0�����r�f2��S�jO���L3M6l�
�6:� ����6���V�X�*I�����[�)�٣Y�e�� �;0n=��}��
�˘6,<�]�;b��H�2��ᦦ�ݫ�o<?�Vg.���q��2��������a蘆�(��8���1��jzU��s��(�ɅI�샎�8[��G�Ml������E[2!%� Oi�4L�������6/�T��*bB@mSV����Z�C�]#.Z��%�Mf�3��f�V�����x�����Y�s!]�8M����IM^$���J,$�7��B���@%%[��屢B�>?[�G�Qh>u��=�ǎr���do�V�]{j�GI��eIQ�Nŷ�y�(�0��Њ(�v��\,oބ��\�͛�j�6��Ua����O�����X�İ��!�|�w�|l��(^�ѷ_�AENv���P^��7��'&����#�^.��g�n���ڿc2~������ssFZ���6}�ٻ�_��I���ZgQA�3�Q������� l���>T/�t��E�[չ-m����[pw'�܃���{�!@�@pw����q�y���;_������^ݏt�Z;m�;a�12*2p$Nc&UsD�U�(�7�U*#1�!�L���4]�����u��Ni����i��|���z<{��i9��BD�;�Y1g$/?d��vՈ<Aa�R�@p��_�}���j0�L�p�o�jHz�w�����1��y�Q�͢���D�2�����յ�+�ʵ,3y=@�K �d��e��gr�ou�	���|��T޹Tl���-����2ڮ�U��-�I�y h��;��P�6z�7�۫�&���D�6��r��q����E~�~ 7qf9�KL
&}�E�R��y���~;����G�>�E?�0�]�����P��O�	�� �$$[��}}	B+���qA/��{E���^�*#ėA���B*:lx��(�_�F�d�s ����c�xl]�P���io�o�4��V�/���\�����Y)�ə�Ѧ����t�|�o�p���8����ww=��Y�pih���&��Q#}����ͻz(;��3�N����m~�����\˧�u�2��a��v��h����4������������*�z·.�������6C4��r~�ٙcF<�����>��Q^���������1���Z��J�_��
hfqq��
���Q��Y-n�x�K@4�0w~�r0�_��`��#_d)�/�$�"���ԩe�<�������wcHnW�2)*
bx�|����$ͳ����n(���Q_z��������Y~M�e_�����(?�ď���e=P���q��:�j4�J��F�k_*dEiZ�Zx}(��16p.�������>�{��ys���V��蔊������S��&�e�7����Y<���kO��zB���V-���>���Zۥ:O��=�̊����"��0㋓C4��h8���fL{G\L�|5	'��wg�yuV�ajV���7<ϥ�-��+�<���k4�6G��^����p��+���S�f����,տ;Y;�,��叿[@�ؤ$�
�n�ё����pws7�~��@��8�K�3�X�ޢNۢ��X�w�)>x�Riy6�=5H�n�g�[o�@����Ϣ���H���hW��Z��yҍ��E�Ҧ-�*�㨭��y2�%voTQr���@�/���������0�.���Ɵ�=�c�]I��<d�(����ot<�ȷ�&��i���i��U�����A�+P�f=æ��<17�&z;��4��NFה�>Ac�vqqY���Y����+���/,����8���f}��R8~�)��+%����A�Ǉ){�C��24?�@�;!�#+G�}"�K���nn�����J�VTE�~!�h�y5t�̊l�R�ܳ?5�c�A�#`�l�N03|���W����x�5�{f�|�R�-/ûr�T��:{`k����nV����0���i���Z����g�r��|�c�&S��Y����}�2?��T���v��*���m�W��l-L� d4�V�x�ɛ,��3`\0k��?;B��оA�%�����
����&Q��X�P2�mW%אc+�������D�^]t����5���`�;�@�55�f#�꽽c�s�J%�ޖ��}�~o�!R��wO���������ʱ�,o$C?W�3�'��;=|�U�-��	��Ax��/&�Ҋ����?8n�iDQ�u�neU/������
+���g��'*#% uAk�ŗ0�D��؇�=����ڷ;�FoMF\o�&���@�ΡuG !��~6Uΰa��)o(���mΝr��C�0�d�����S<_�!�w�ր�g�ׇ�����|$x\��nǻԍ�7?H��ME��G7�'��0C%��w[G,̻���OOz��I�إRf��pN⏱�i9hRh[���DP�~MިQ��$k,,,b
N���g�>�^�飯u����z���9Y�yQ����m��ң�fܻ�Q_\�v��N���f�=�ӕ�l[n`�0�+�c=쿅���H�qֻ��iF��z��`����̂^�$]`Z��!��{Hv��b)�4�HB��>�ZS|�8ĄX���Yt������4�i4�.-����u<�j�1�	t'�$[q��l���e���-�i,�5��~+)���	SXR�a��[<-^�E"��ǹ}����vy����ְ�ŵ0����7��������`oc3&Sި~�B�S�GWR��9�P���R��N����*��
��/�C�orB�^�i���ͪ��/.���jp0ؓ����f����ʝ�������Nly:�+����6�.C,���!��/S�O�O���N�쒩k�Pϭ���&�����7�8cq�����O��	��e�Y�?D�ġ�׽Z}ܪL��زZ���7���+���Q���B3�?�������@當���/�4����͔�U�>VP[Gſ�`�ǣ��~�IOe��/,oܤr�x����	��g���}�h��YKh(B�:��l�Kr����+��1����.�\��� ½���s��#Hߛ �um�O�)&�R#���b��[f!��/[�q�?5H�C#��4u����^t��t�<�ݯr���k�IN9}�W������P�@;|��a�������b�����f�X	KD��t�e5d������),�}���{���^B��xm�~�;X���2�.�Է���}�^���>|@燎N���H`=}Hspb�����I$\�*�����1>}T-���ҵ �`8�mW�n{���7�x67T^�7��o�A��%���zx��� ��CU9Е��s�i�qK�V��}F�F�[��� ^�̏o�D]�����c���k7�	h�_�(�}�p��o+����>�_�>@�q-Np4h(���A��?��?���lc��Þ�ã�AtM�@��w�fq��� �M|FW�@�E-7�A*��������#������$��ߨ��%�6.����&�C�����q��V�7�6s�3ݠ��F��I����[o"E���fu�;�UM�b���ʅ��M�=Z��S(Ivvj���É䛛�F3j��Ń/��
%���{G�IG(����e�l��N�-Q��dC���]���D���H�,\V�앫{/����W�ᨨ�S��/FN�=�s�Lt��s;/��<�NyiaQ�ِ��퐪��AW=�F#�:�S+1EW4,�M�y�qz�$m��0��ϐ��=��RR��iB�o���>_s��X��R��[?�no�|���T��:�F��q�p
ͪ%Ϸͭͅ5/xx�<p447���OS��S�^y.��b��k�H���j_CB�������d�\�o��n�~�Ct�t��Ġ���?O�Q�\�#I��YX�=���/@�ا����p���R}����s��ۦ��	�$i�P����][�/F�=���p\o(��Y��5����jUs�������j�����q�΋����G�����M��%�nT�"ʁ�`�q�.�L^/(ڸ�T+;W��c1""b�I�(-f�*(T�NA��J�y�s{��G�a��J(<b�{�f�k�K[�!jB&*2�ElA�@�^�E��&zZ�i�A B��:�U W�-��l�f6����P�.UU՟mm�((B�)����X�>|�F��^��W
D=S|,_���'�E)�#2�t2��vf\@��øJ{Hc{�.v��L8-%U��Yc7¾L8�hU�A�9@ߟ�ȯ����2��uS��,z�M�oư?�JW�	ڀ�$���q�~I���@���@�+���`���~#��^��`,�����v9(�l4�![k1��%�H[��Y_	4�/8�S.�z8��T����M+·���.v�p���7�gZ�9��v]�RR]�V�Б%�G�~:���Pһ�X��p�~)�hjJ����
o��+�e͍r��Lj�OhU�w�:
a̰�/�������j�o��R9�~��w������I��a��Ì�ԏ/�	����KsO��EiX�&lk���w؏=�j��1�9�Ne�W�gq�3��b����Ǵ�1�䕥cb*(!|�MMwT pf���޽]��SYPF�[�z�G�c�Ϩ}��P\�{�s'�'����a8�����V�f�3Lt�8��ܵ5�}!n�(��9Vg��WK娱+�G�aq@E95���m�e�|ϲ������ŧ���@j^꘰��ŷ+�5���3oF�7��-7��B�@��E$A~�%���oH�tҺ�c
b[�L�-��p������bm�?����n/�XZ�=|���?n��T��_���݋�M�1�[����B��(���%d̋S��3aeu@��
۾��z��1�P�L�tn�Zda����\^Ӥ�h%��l9�v��1��w�����CE��N���f�a���}_��?�/��+�}6�/�[[F��/Rt��:І$��56�UU��.��˫r��}�����'��5��\Њ���LM6!���a-#]��t�í*	"B*��Ri�=;�ߝG�fS'>�*����M��o'Z��HEwTTɴ羾Y��2D���L��ڝ��ly����ޢ���'��Fr�쀰�F.c�!�A�ꮭb� 9�g~����`0&��������G+t��]a6ߕ����p�w��0f�@ɬ�����P%��i�NNm|��G�������Tt����8$�{�n߽6�A�sIe%Z0,*?�DP��������^���}�p��;L��'8�LrC��+Hpl/�?Mœ���lH�ԙ}Vth����s�l0����z�^���λI��5<!тT�����褚�
r�u��H�z8�_�y���Cr�KX�P���l?�����0S/���-�2]^\�B���<�ό%%U�E
٢gUƼY���	�͛�_vs��3�B�Y�	
?��;��lƤ �$�6�X/̟�� ee��U��\��X�����&��$�����]���-m"8X3����� ������ ~�:V�i�#S�6>+xz[Eu����F5a���}��1��|�I�������1�m���B�N�F�Ht��M��Ҭ���3���Z�������ć�{�qW�#�[���i�,U�>�����vߋ3·�/�F�\\jj�N�����۴��M��e:�*��u�K9^.���/?>Ѫ<�ƩW�f��$J��4�p/2�����?��!z����qx�v��u���.��!z;� ��\S�ǐA�vv��2��4���ʭ��Bmrg
za�
^��c�b�׎2�����y9�%w�!I�·�F��G����O����i�p�s�r����ʭcD�Jͭrq�Kڅ2H�HӁUY��wt���]]^���O̻�|��v���9׃N���_�%Β�Ia�g����.�.12^�"�}I�<��ڈ@���dy�l�.4yT���e�0bt#��Vܱv[���N������6m쓸�Lh@��z��_�5�:�(�۸�D%���Q��<��T�B���nFJZNALӃj��q,k�ǳC���<+g�y��y$gG�����gf�e�NÌ��fs��"fw�\w��D�=��|�.�X~ofe&�4�n�½��us0�+{Fd�WX����^ٟ��@��x| ����'Q%�=&��D��4�Ͼj
{�9"���3�˫��:H'G�+}��T���w�q��X�7����'����t�	�B}��&�<�{!srkJ�S�Sal�
=�4<��ٍ�wf`a	_
���&�K�@}K怼�(Z(`��nh�9�f˭J:dȲ46-�F�6X������__:-�m��Ԩ�����z��AȌ���64Q2�ܬ�ح'�}�挟�9=tW-E�/�7��u�QY�ʹ�6Q�v)BOO��y�����i�ԗ�3��t�����k�����H�b�Y�����+��Q_pDs��q�����v)Il��M��mV�K,1�)��7��xɞ�#�Z}��'������F��?��L%ok��W�U蓋K�ba�
9����MpK�������φ8��ܒ���:��%?v���-3����_�iJ8 ���ԍ�[&b��j�)i�X�Q_�q�ZҶ7#{�J�mxo�r�z�,4�B�ȏA���fN�F��� *�1k�����E�޺���m=�2-GǪ�����W����\GNV�/��e!r3;U�gӏy�A�/�e$}և:��@�	�!�/��w$��KAן�&v_� &�FZl����\���/���h'�9g?��f:'B;�h����S�*�}-�T9�4 ����zBqш��\� }�'���q�K��NP8C�<\F��,���Ǝ��w���^:�:�Ƌ��C�!���L�CC��K,�	�R�N�!F�"a�U�h��-�6&�ơ�s��v�l�����Mo��0�s�=,�_%�B�|�ڋ즒X"���MkUM�4H��^�i��8�<lZ�>�-�u�L&"bI�=ƷoU6�^6���
����s�.�Ņ�94У(�s���ike��o�C�⹢o�C�
�>�F��i��;;H ����S��5������A����4�3����yH1W����:�����\�"C{�&D��BB@���b��_ŗ��|���v����G�1���S���|6�\s� Ԉ�����V����0
&��A��5��+�Ze�!��!�L�E��Gmh�.e�,4���Q9
����cyb��幑S_��3���D��+uf��d+..�@Xy���'@�hA��<���_��={@	��-��w�ǋ���"8:v����KWRu˃�����YzxPt������mW�e��~i+�Iȏ����g�����E���\p@��@G��a�Ј�757�ٕM�|YZ^�9;��#¢#��&V06695��β����,R�;��,�6�j\��̿=��5l7����X�`3�8���j�L��-���I���Q�(�q�;��P��~��'���\h�V 6� $E"��NPr��Gpb�V:����Wv��
>Y���񗹾"E��I����7R��!�v~�q,�p,e�5� �~D0�[*t	M��G����6���2����ĺ6�
E�4��bɼ+?9�夰��>�O�
�/ϼ��Ǜ��{
�T9̨?(C���-�n�B!�o��byW`�!��q�������Y���X��|YJ��ߐV���#ַo�F��ٖ��͆��Pbc�bm��50q�E��DѴ֪��[��ۭ��~K�I���1%w�V�bJ��z�rX��sC�K�:�S(M���)eHBv>l�������̇\�J�Ùǈ��������/���d]	������� |Z������	G=HS)��������
C� *�F��=��kB����%DT������ ���y[V�����q
w\I���3��N�E�֌fj:y���$�?�R~~����/Ed�K("ʘsM>Q�L���_��½6�}���P.�"����|� ̔۾d��ZEu�A�����>˔�bTW�}!y�c4LJ��>�v���uw���t��(�����a�����OW ��<s������� �˱�A|�d����V��W�C���f,S���W��˩����z�P���B!�fM��:�ȷXJ�4^�ˏ�?\�D�X�8�ȅ���w�@�H��� 4S�n��8��awa��ȵ��_nS\��6�꼉q��h�ؒ/ޤkr�)�S��P���{��껖$R��PJZ_��#v`r��&D�?H��uې�
rO�{��ז��_f&�`����B��ͤ�X��RG	�#8������MM�q���i;SZ�I��M��W0I���Õ���O���7p��}�����D'/�Ϧ��״X�Ɣ��\�������(�s�|\�Qݥ�����U&1U*?;BCA��L���ೀ(�@0g�`��0��_����=�x�Ilѳ��,-�L��6���H��������Q5����*�_�����|�E]�p��P4�3p��t"o��d
���~��Exk�K�n����O|�쁽�ݰ&�=��xg�P�R���yB�B��B��j�:����&�/%�� ��L/H1upӺ=PV�IF�%���tu�W�trɪu����X�i�,Tvc�x�N�����$��˨c�\\G(!_�^Y[���h�x��Y`����PYY�܅@}tR9P�P$6ǣ�GdF����o�s���"�ؘ_]}����z���H�-ޚ��$z��N��H��̈�X��L�獻wRݐ#��n���p;t�_!�@;1�d�2�k:��@.��YД&fVx!���'�L��M�A�&�2��'F�վ>nTB%�?SƫQ[Ql[����m)�p�y�k������$'�|z�w
F�p��,�x����q�LdJ2O :���V�x�I�c8v��L� ���FGjܾ�1�;AOQ�w�s���-��<X�O��st����v��1������e��#��$�8�wn�w5O�Y��n�qr�m*8	�H�N+l{FhI�+l�;&��Nhi!���3����=d�5Y��A�ǰ�z���Yo�h�8�aII��7uu��w)=���)n����y}$X�-"!�K`�3�vww�n��`�}z��W��𰄃C儥f�u�f�q(O�����ȡ���%�����>	��/��u��:��"�D�{�8Ss�E3�8**jJ>&d�XQF����AA�G{a����K����SߌB�B9�ʶ߉h�ec�E"��!��p��7�!����J)�(,�C&�ݙ���sxK���}Ci���𿢠**�4�x]��IM>�[��w|5���]ѱ	�m�##����rϚ�b�d��}
�&�h��p��Th���A簏�2j�}����#0Ӣ�_*P��UI��=�ț�4�_�dQ#����$3����}�!,8I���?��hK��^�X	�ǹɃrL�n�Px9}�'XQ�*x�٥\D� `q�� ��2a�i!9o}�W�4���R��{�1m`No�mv��.�Z9��A9���_P.Z�ל�c��F	�<R�Z�`$��1���U���`եcn>�yl��!		�{J��d$�	 �M�Z	����-w�~�;//�+���U�����TWwu�p���cuec�Z�G#߀�?����@�0o����ޮָ�(���{v���N�ċ1�! ���}^ij�5�vLH�'=�_�K��i��U!�滝��		�2Uf�B3�x �
�h�fy��`-�>�	0����"6�fw��ۅJ/h��^:�i���G/Ι���_���z+�o�	�������}���1�
�|f��A��!7�,���W����J�켎a�$Z����% ?<��ލ��
���ı/}k"q4!�!���&g�NiE@��cTp�{��}�w���U#w�"Ê��_�\}�4�|�*}v��/��7�fAJ���������\��xuo��M;P��%lO�p��N���W��]�Û��$"^��WWNUF�Dr�>���&	���7t@)e���{tn��)�D��2G��y���R�=N��	K�� ����	٥uq]��������f�����9����T�����q�c���h�� ��}��@EU����HV��B?�v�v6�7
@Å��Ă�E#R0�[+�����u!���J��cQFm	jK]�m�s[��d��Պ.ڥ��G�H!�:�"Q�}��ޱ_6X���I�(�S�ߌ-�x�;�'b��;�h��8��݄| �L[G����}]��5��ҟI�j;��{3���=´\�]r�S�����Vu�Ϧ�2��}j�<�� ��{�7�������l��0Nn<��nWBL�Xj M��c�?�b��̴��Ey�)���hM�j��)��>=�����#�IÈ)��R�@c0�{����q�qȪ7�@| �\��
��9�![���͇N-w$�Yøiw4��E.�F�z�>��Q
�匐�[���6M�LC7�$ֵ��Ǽ��Y���t���>nNa�*�j�j�>ŲC
��Y#j����ww!����q]�=���>�����X-�o#7�}����^0�4D��\#�\]�����  �QZ/cg���ܧ)���MUO:{?�t���K�����`7 /+��F�G=��<$��#y/�4��i��=-�7��.cx���aN]���6g����r��������!���2s��WX{X�O^�_i1([7v��+Q�4�64�O��e�&����t��N��f����\]�;P��ɹ�{�+��,ֶD/W(î4���������}������O�o��H2�A������W��I���՞���,R߀u_1']�l/C��?������zt'ʶ����'?e=����l	!�u���I��x�bxB�b��Oe%ϖ�I2	�u�G߸V���o-��6�8o��?a�,��i��VA�>���7B%z�M7}�i�]wT�X�M��3��������ӮE��²��y�����R�l���_҇zU'Z��&k�o�E�Oc���(-S�QPP W��B����5'|�~���;#o�T����?��v
�����qf��ʹf�$���Dߣ�{�*#!�D����Y��o������fI��b��!�O�,���J��L�#/������U�����$Lz�_������˃'��MË4���;�ԇ�s�Ԑ��JW�8��>v�U�a�Y䅕,%"g;z\:�2Ps��=��9}s?fy�[�`v�H���LQ=6/nnL�I0~58>.���<Q�@�A��nݓ�+!�'�����H� c����"� ��a��/''7�/2�c&c��?B�zS��x�&7c��k�7��=�fs\U�۠�υ��h������Zm&�R���a����iɊ�[�o�M��b�����7}�-0bP?gY �d���h�z��Y��L!��"�e#����:�����~�xZG:�E]�=�z�6�,��e �/0!T:��ΚL!	�����$k9�t`7Da ������a'�y̸.]@ً�s/�
�|�5����q�4�y�&��Z�pw���*H�p!%M�����H��C�,PK�[�ƀ;�������F���?�Ĕ��ŵ�Y*�k��lHU��up`�v��o~�7�A�4��o�H-�$Mg6ҡ�cG|�<�(d3�}�\��0�����4
N�\�IZ(#����n��.�d���ǯx��"HU�ڟ����ڣ�%��8;d >lc5T�Xl�@J���G����ڨ9��e<~�`�:��"feE�K�J)�(��/��F��9}�[�J���*�"2���>�IPTU4��F��ߝ;M��'����[��,�t�y��q�x�/��\\%ݹ��ף�@�Eĝ��0X|�!\��:wrY=��<��Kж�`�O㙪cW~�����(F:h���О�+����fs�1YK���@�WE�U������m���KO�c�]��X ɜ�zD�y�r����F�\��$�u7"//���Vs������Y��ь�M��*��sc���]�k�4a���h0~��n,�[��<�:=��@<.?rFr6z[>�n����������m<Id� �T��<_S�A����~�ɅF$��-�j졒Ä�&8�>�o��������v�}�7�~"�s��i������e�kN�\�tO�j񩂘��M��+bj����}�Xҙ�F���#/��CI����v��7��Rx�8~+Xo���zz��zG�.yV���C��J��Aj�i�QEh��p�0������=i|/���J�S��艚�G�>�۶D�;/Rh�"�0��/��6.'�je�%)Ѝ��]�"��յŦ����?A(�����hm��>?2c�F�ZxH���H����.|A-�)�� P�b���=?���"m�H�  C�"�?�hD��g�V����^)3�?��3\ɠ�<S���㗥��_Q*���.�o���B�����[��;�muAV��\�/��G9A�%蜰��TT�w������؜�Wٜ�(蟉��^}7N�"�O�Z$�7G��XN�;DGt��}_����1+x�3G$���r��h��c�U�%o���X:�$�h�ء;3.�P��qq�L�(�Τf\,���JM>Y�TY��rW)�E���r�~��A�]�Y
��M�����(U����h�.�u/�Asƌ�QD�j��9����&�:�M8�����}�^5@�\�m���%(0 ��	qq/�����S��M��	m<]>ͫ6G�"�@�s�X�T��0�+^d4MDD|1Q[4��c����.}����C�{[����Q0�hQ�o��p�7�FU�.*��5�xkm��S}hQHPMe����6�+�;C��YGʎ)��،�(l�kd
6�5 q6XlASgf.V���A�Z/� �����I���$ޥ��ƍ�$%��v�u�4�y���ōԹճ��
�*�x������w�J�;`��v@V����hG��Y/��Etŭ�R���0��'(�'��b.ϣ^EW�5����p���
6�����ېo���紙��y��)��+�G�
�d�ߣ�fff:��u ������� �y��Gy��iXLg�؏=���E��=i�Hp�N�� �v������%��������f|җ}�wG Ř+.s�#�J�.�AQġ�f8i� omYkG�[���kk復��o+�GdK4�K_M��'�J�:�.:Ma�V���~��=}i� �l}B
3ܵ�׵�B#�PGt?�k7Ӕ�!�ܹt�IY8���R��{�_��YQz�
�R�M��c�V�|���S�ϓ��K��Z =P]�����˓����d2��|��ٯ���k>�$�0���@4@Sew�Mh�7�S���z 
o���2�{����wV�L' �����}��ɭ�g����u��@đ�uZ���z�qB!e�jSY&�IMK��HX^� ���.�#|��e3�A�R>\�4Uk t:��ߎV��+���̅�;��*�����X���rF��&d?G,rˍ��XĂ�J���,2gG��d(�s֮��R��W?��@�AF,�����x�ú�_���`�TY{�d@���Bs�25@��v!yCxy�$�V1}Xi�_�_�����Mi3'v����Ow��Nw���婢�� �E`�k2v�x��g��U�ai��3# xx��:�M��a�t���4LLTi��`�j�QYP�|ca�j�V����2cR���	�B⓺HR1��}�'w��PV����t��	��u��QV&<�(t�mĖg 6w"�jSt��-|��3!ܞ*TE�ITv�@�Ż�#
|3[�u���͉BQwuMMI�j���������,.1�X��8L������^v�&`���0c�Μ.�#u8�N^�Yz��6���y����x9bk'�4G~���u�w�X�%2쑿�>��V-/��$Y���gI.�����Ӷ�yL�+�`kk���Am��)o��c�&����1��YYL�Kɩ'(��Zt����y�n�b��߼=d5c���J��x�U�q�4@�H}���p� y��z���1��-]���d?Z[�l%I?���7�C���v����G�xƀ�܋�'�"�L��N���-ճ2i7;U� ��8I8��|�l�]�ꆝ�	���:�E;����*x������*ǻP�;g�@�.���R�m��w��m�v�'��#����l�y�2؆߷�.o�:��|g�f8�:G�||^�W.�����%����?��BjS,%�+��|eq0C�H�N��6�.S��M����r	���j���d��QECr�'J�fy�+D�r�+<Ê: �g����-���>p����s�~�Ji�|�ϝ&Yh���Q/2��5b��k�Tf�Zx]�S���&l���Y�����q|m.>^�����g�čMڜ����?'-^��@��l�]�6n�,����a�?m��%|hi�2�����X��½/����48D{�J	/���iI'ww�=С��}�x~~q�ĝ~���]},�O����G1���oC��^\�J���׷�����& �S��G2y.��r�k��o�����I았�~�h�w��+.�*�[�,h[�H��i*U��``��]�?�&H ����i�݃N
��r�m-f��������5DX�J��o�l2�^��^�5�Z�y��+Rt�m�[33�2�`ly�z������cy�$]M&>�F�W4X8�h2��C|�򅍕٩iŨ����g����^Mќ|���/�4�4�������M��¿�G��ص���F��@����oX���^�<܁�7��BH~�ϷW��'\oz�!��?⛊U�3yW�� ��W���E��p�
Qk��C<´l���9��\�E��g�pϤ��0�\�C�Pݠ>w���WU-r.p�neyy�,��~�	�ଅFF�6�7�m�`�o�8Lr
z�C���o�P(q3}��~�ɵ��<vy��.�b�oe�#�&{�7�b�����M��Z[}7vO)]���/�>-�eLz�5�qG���N���G���}���ŲH�.��;{��%Ь�O��*��R��%���1�	3(>�#qm�H-ߠ�ҹ�ry��[t�L�'�|ƯcqhZ.,��Xָ����'�������l�ڮr:ԧg�`�_Q�P��G(�L+3w�RV=��o�9�J���֒����<�`�c�`�G~*�������z�J���	��F�t ?��R�~����:���@)�`i�������ۮ���*�Y�u�,���_<<<�2�V��?\^�<���K�#�#�O�y�A������,��T�	��>U]Nc*Y3�8�s�08��\i$C��#�P0�K�2{���t��N���&�#994�!+L��ѵ�:���}�n�a�i�J>����}�:�V�۳q�I�¯~����$gB��~�'��%q�K�+��vkw�ҋ��� Da�����_A��H��W Q�����~d�>Mb�%�ݝ��t�H�b�гl]#>ص��i:���a�it��GC�i{z�?�-���MP�-�t��_���
�D�:9�C�r���,�#��C�ne7iȏ<�^�&`WMvƁ�e���i�����K��ٵ�<G��nK�Q��g.�I��p�cz����ǚ���S��S�`ȳ��7v�NDp>%I:7�,J��}[`��z�
���ڷiJ�A���E��o*�ʜ�`"�wȒq��-��"���l,�����˴��D���|��]��iH�KJ�8�I߯`iN��P�&��r�~�W�k���2>�.�ܪ�i@�aT�ɞ)Tn�vd�W�j	?�i�I���t|�]����d�A�b��O]0���y�}吲��/ʛ׎#�iL�V�4[P������Z�{��@�	��`���7�t
�v�s��}SW3B��p2��Sz�;A[���'��T���W��=fЩc���S[�U�E���F����x�1�J1�k\r/וOഹ3���F�^��ɿs�;\:��	�b� tt�@i�H<T��"i]цF�f!� ���%ݘڌ��Ln���{@�v ~R��qyg��YP����Vn8	?rˏ��8PĚ��V?q���< (�Xc2 ���RH�?R�P"D��D���͹˨̠.3je���b�qy�MKKK�H�JSEܶ�Q�p,e��"<ω%�E�VN;�zSy�Hanp,L�C��	b�X�𩓻�u�r��@4 �sU��s7�sa�����A����}X��i�.Pmt[W]0�uMN2G/W � ����:lY�uywSzs�Dh�>?�p�� f�������6'�OD	�vx�k�ڙ�q,�{7`����!P5� y۪����]�M0S�����Ki���W���K	44���G�P����jTo�e��U�>F� Mf�����9���X�1ø߄��ZG��v�mܟI������6�NP������&���D�)1q�����>K���ۛ��\�?�����Ql?�"���:O�O��ӟ�����z}}}�aϷ�����L�oKY*���6<�>>Җȅ��R�25!+����+����i0���MCL!��{�9�GB1KE�ROa���lz7�'ů�~5���Hw�+C/�G5I:C��<�g�qq���<�@za>���E�:QG32W��vrvN��dt�wS�O������*Ǹ���\K�Q����7'd�P0��� �9����F�ń�������>p�D�׸v��|z���)��FT	�D�s��D=�v!�����P�"�umg�z��1P��1���>^&rWQ�"AU{%�s��d)p��r�}�ad�/d���3���sr�����L�tM�� �~:y���o���#E3	nKh^�'�c�LM��[P�=�����	�}�̈���z�i�-��Qr_�LE7(�>OQm����|������F:v�S�{J:�������Z�X��Lͱ.2^KCGVą��)�lVh�V֎�����z����k��	���	��!��<@pwww��݃�;|C����_E5U3sz���ڽ�ilj�P+l��+{H����f���~)���خs����a�W=�Ԥr%��Ĵ�jňB�sg����W�Z������Y\zm�����~�Z��{�h��.�~��n��U���(�1�K�Ҽ;u�- �o��l~������j�mi/�uJ۵O�v�R�U@i�v�)2x|m���<n��"����ݣ8F���U��tE��t��C����P���=� ySܝ��?�$&�Ua���6�"(k��QI�B�4��ŭcg�C�ϡ��v������G��WYZZ�}vϙf�/����c�M�MGK��a���V����3�\���������Îo���  W��{2�'���$���+���[?�y;,�=�7�	��#G��S;����К�߱��@ݜ.�7�l	2�����c��0b�I!o�S�GYC���ۆfIЃ9^��
D'�����ZY�'<�`�N]_�|�DO�e����!q]Ά�;�+���1�����څI���{h�;��;ԓ���\{�//2օ��l��z��IX�����؉ѫ��2= L	'��w��|��`&;��$1�q��^�lJs<�|�qt�"�.b�����t>�}�ւ�������[[2�I��L��2 @��q������
�8��=
�]=h<�I�w��V���;�pr2��`}a���\.v�\D�����Z����<���Ne�ѯ��:pI�/���6�]�CX'�B�2^��������c8�v�	��\�z}�U��b�v�}�?���V��qo��b�(8�}��B�Z^N���'^�h2���齆�Ζ�X�9�:Ib"���^�t��򃘇0�A��G��b�93����U���Ȟ�󉗍 Y=珙f~zЃ�:���T�fQ���q���as������l�K��n~g`g��~4�mm�*X�J�˙�U�Շ�����~�_��Ha�&W�]z�f�O�9Pt?���];Rd��%8_b���>=>ޖ�`�/#�d��Ru��v?|�7
�N:�lp�ϙ��v���1U=�]d.d��bߙ'l�dlXtu�X�w��m��ϵ@�vȪ%'5����W�{�����
�����zit_ �cߴ�m�9G��5��^����"o���~g��7p����$_��S^�.�� L[ʍ��ax�hȯ
�@�*Q�I7!v���f#W3W��䎰Z����$&�g���N�N�.�M���LF�Bч�h�|I���OL�eڞ���T,,h���Q11)�i��~z�!�-\:��R}.����JS�o|^�	���֏zS������&ѿ����,��/94P�u�I_�O\��`���4YA;���#�FU��0�z>�0$�C~6�S�sGRCP���p���y�}rH*aOk�ls���'�z��V�(+���U���h�����71Up0��D`{#�U����P>=e��/��GAd4e͖N>6f�|��=�Ŝ>�G9>� ]��f��Dv�K�ku3aYz������e��g�]; EƋW����Jd<�)�Ҿ�z�6��1����@�c�4�u"��������ăC 9��GO򇧶�nr�v98%��3;���̯��*i�Ye�����r8Jӳ{ϓ~Oc2�?��F(���y<� <�3��ЙV0c�v��j �~�@�boΞ�Q�i�ޱ�|cp��nx`C6�(��:�o z��Aۿ�s�w�u�V X�{���m|X�F-��u���+П@�n3b�
8Ī�d��jM�5�����/j��.>���`\��&.}�����_[?�+C�x뢭���_��dW3�ٙ'S~�dԗ�b�ɼ5�*k{g�FQ8������o���K���������A=�������@�/�)��������9
8��Ad��F�����-'��;�-�?�������ߙ�<Uc�fָwp͗����ΐ��]2]u�v���up㇜`v�CU.#���u��{����ߘ3ӮWq�4�4��'��
&�����*���G2#.^J�I�J|��Y�I�+�Y`zf+��|���Ǩ���=^,̚v�GrW�����Sr�AR#�J�'�V�J�c$	�S]e�j��f-��3��T�ޜs�o6�&U�H�w1,`_9�2������ڞ$K]�:#��u��1�3/�$Aϫk�����$(

�w2'A�����������a�C$"�0t��yx3�g�,֞�:^�0q�����l��T١M��`�2��u[v�Q�  w�G9�s���
�ݫ�8���Mz����|�i퍤��x�Bqay�1�6�Æ/����y��Eq��|lTt�B��!Sf�n��6��7|Vi��qS��@-
2�bH��$��u�����n�h��>|ė�TV7�������b��`�v#�J؍�*5jV��߁�X�fe}���X�0**8����'-��hMmZ�ݙ����xh�?�R������+�9ɸfqz�ҧ��Jʡr�Ը��2���j��������g@Iu?��MHT�YOm=?J�eQC�Y},�7��u�I�#	�U���	���ĞN��郠��xJ����4t��*�^2�*r���}�{_���եs��%��I�'��(�����(j"�������@�n��@U�V��9Lz�zyQo-�x[;<զF��:�9�l��76:fl6�]���ӡ^XF����G���P��x��0�:����1�[���Y�)?:)�J5h�޷�MH8�s������I�5o����spl���H�6�7�iq�&(�*��9#����XKq���q^�gp�J/��u>9�}��x)8�NkEY��JGp��ۻ��0s7h4e:����tb�L�:��rEz�Hjd�k(m{D��<�ô��#��z},���26�����#���ˀ��s�����6�����I�v��	�!��K��G��V�t�o|�\֭/��*�ăQF&שۼD�{�;^ek�O�<X�Ү{����8����4�!�����zqH;�<�+��^Fd��	fL3H�= �q<�a�╦Y�����J
zj3��4O�si���㳍W2b�y`�-�d���:̶��X���}��S��O�Q~�K�5�(����	@�Q�q���4����"��A�v ����j��x���ec�W:A���G8v!?Eab�ص����@��šc>ޡ�ה���8��N�W���t!��D �{�M����$ւrV`��#�A�E��K��W��C���`ڕ=x�|�EI�T4��!��O: ����Z���K��eSx�4-O��$N�6LK1x�iԪo�W빽��݁�W�
���=��f�lRw^��}�D�y��u*w���Ι~�.'�2��N�ḷٖQ}z��<��Z���Z���7U'���3x^����Φ̝^�T��#O}�Aɏ��	�on�9YA��Z(��E:�ߙ����L��\�&F�0&���a&���r�A�yÊ�{{�'�5`�X;LԖF.lN`��9$❦f�ɺ�A�m�S�m�7��N��^~=ϔ�N�a9.��0g��i�z����D�l)��ۄ?%��+��j�����t�>a�Z/7�Ě���=���u�}�����W�I���1���;=C�O;a������c#<�����m�C��g2�qL������<=�	G������/�����o�eh��&i_g<+n_N^!�j��Z�$0�|��/���KR�ɹ��������b_�S���4!���s�c
v\w0?f~[�ҳ��PV23k���7F�[7��U=�ot�Ͻ���z����n�d���v�_t�ۦ2"bq7�\7oe�b�{�xk2�����V�cg;��#�[_C^UO�U*ԓ�j��e����a�賟�j�1G5��5�f��g�����oAA�L�*����=�'VsN���z7����_ݽ��սY;�e���M�{ ,�.��Z�^��~��3LaF�=�!,)���$h�T.�+��3�o�u��3��(�ԫ��9�ހOO�l��/���c3b�F��.�ݵN]D�V�t�jɾB�v�l�Pz9�i F݂b4E�;�3&��u�f����)qE~�XU2P,���
K"5�c�}�#� �6H��ݳtp�`E�x)5"��l���r0r�ڪ�$A����2��I^��Q�CpT&�:_Rv�Uv?o��O����(c�0s��p�J0"L����F3�*���e��r���LɆj�.��V��OhhZ@�H�E�î�>e6vL�4އ��J���Q"��wrr8sؓQ/Z@�G[��>͉�H<{�ФP�3� �&rc�8s\�2�������4_�����Mo���"�C�T�[iNMy�u�yB��]�u��MP[��.��(�	-ma��?8rx#d}�OE��|yޝ��T��Bm���ɋx��B�?�{�����������C�1^�^��s��n���߸}�<m���S�`���a\'�C<>�V|2[f��*9�l���D�=ͷz�(�͉�,���Oi��y���V�g֤d��{������"�7t�W2����C�qz��ή��W��%�U�E޷D���XX&o�/�!
�~��۰Rr�۲�����<�j�_"�����+D響�Wr�!�g�Z����Yպd1��W'c(ZP�N:��R�9�>4���5g�--�ƥX�4u4��h��P���V�#j��Z&��q�� /w��}vw ?�=��y ?_��s�h�r��M�s�9�FҩK蟟��nv���9��9�`H��1�܅J[�P*�2�n�4RG����p��3cv=H��7kǧ�x�^��IA��|�0)���,nN��V�E+����Ց�(��g�'A�J��M����A��u�}�>p鞾�ʥgg��P��z�
�������o�+9����t�����2$�<n�剻�lhpEH���������0��z%܇*�uTZ�Xb��HP�39ߎ���h�{y�(��ܽ�}��PUY�<׳��<����e�� ���S�:3K�ȵz~\iݍ�����L�_��b'`��b�*z��ozͥ�6�`�%B)�0gŢ~g���U�xڡ)5��J���m� �AG����pL�1��
�ݯ��S�;��Ԕ�CV=V2�ζW�3�f4������cz=�}H[~�Z��w�tfK��Q]��_ע27�������e.)��?�J�b�NS@��̔��x�뵚�:�j=`_� ��Ur⨗�]��õZ4
%�?K���`Q���Q���'_KəK��u�#(Y����?W4��OEDh��Oj���C��7|)4�"$j�����T'J�\h��<�Y��)�=�Q:��W�q|	�����N�1Z�e0��"p%=�Bt� ��?�5��)��?�?����[[`5�߱�CE��@&��bg��V�s˦���q�h�o���Gm�mc >�;�s��E��@_����ᩓ5=u����:�ϰ��ӈ^s�mm=�2�U�(�s�zG��u��p�f��#���M��U�b�}ϗ�ڧH@G��Pңe�L�I's��J�����[sl�H�9�-�r��uU'�V8
�R�
���ْ�0��6���`�R�u��T"�^P��7�y;�힤~6��u����\�%V��%�mK0ES�\N	���PI{ؿ8Y�6X��F�&ɨY�� ����y�~���T\�S�U��F��ķ*o�����!�e�1�b�7�e�^V"����zA��g�q~6̘n���H�KcA��JI7"���M�����k�g���,��A�<����ݘ�Y��Ҡ��O�)hO1����Z�So�Z���C��Eh55��Ġ�������@��%�$�[^�o�������S��B��lƧ��{.�ܳ�}l�1��}��
w0���c����-�~&�XPt�=WP������L�����lq4W�o�URV�Yn����/L���|�m���V:ܰ#�.(�O�*�d�;V�'�@�C��e�8�\򻎑�+z�ZKGTɑ����k{B34�﹎JL���}���_-�� &?	B0wV�g\�m�m�"���ڭH�Ci2�J��.�$Q�uAś7t=���^�N/�o���z�mu�U���M�݉�{�p���F�6�������Z��2*�MT�e��r�J�
*�W#�(n��R�^��g�'��������Ο�����! �[tĎՕN��v>t1�+T"��?�~�IJI�>�j��::���Q�|�I����+��@��dmV�n���E&���q���!���OWDJ�W!6����."�?�n��7���Z��@��00����ϒ%Tst���-�
��j�g��&tc��`>u�#oTЂC���M]��~'��2�9V���&��d�T([����a��`����@�����o�.�ے�"oZ�eŭ�K�ʷtst��4���l.^x�T��l�� �F1^����Fe�w^��?�J|�Gn���k��f�NL��0�1p�Q����a=��'<�,Qs1�\@�6�p��&�D�_�"�0���_�Â�G��Y�
���ثkdw�'�c<Q�c�Nsi�)�/�k�{�J��(A7~�~��-˯�mNgv��
�G��z�����h��t��n5Ӂ�O���D���q�$R}�ۦ����k����t)����W��O<!����v�Yn�ѹ��zV�
��4g�r����X�ҵU��q�5��J\$��rs3�Q��^��K4���aGu_%�eS���Q۞̄����|^<��d'IACו��66&�{K�P�b1�e��6�J_��4�p�/�JL�����1JH)� )��:�B �HKU��w���cA7���zE�i���m^��/2�@?�sg��@YQfw�q�<��F ^��̆[O *��*o�Hw�2U/>4 �o��L1������������DӇL��x�w�fV��R��8�Xw���;�Xp6}�8w�}��D�oTr�
ڢ����v��U(40_��Jɼ�q�S)��P�\Ͼ��Hv�i����ÂO��E��g�.�C��f�0�ɪ�w�V˦C2�I'yXR�T3x�O=�����������3�'��%n�pj�d�h��yz�R$�7��� �Wd�roj^�'�;�Z&����e�����q�|=�pպ�	L.jX��r'K�l���r�,��u�����0�T��y�$�2~U��+�m9���ܪ7�OOa��}�7����"Q�4��`��;>�:�"��QK��:5.��/W�_�5������������$9E8���D��1�VG=|Җu�vӉ<[Ƈ8�rk����4��E�>�&!�M�iD	�C�athB���דC��b�t_f�m� X��#�)��rXl.$�6���}�osh����-���%��{B�+����5G|z��yv������qN �)P���r�=�r##Y"�\��)�j�{�Y��x&¹ݛe*�O͎~��wx#HV6ɳ�kv'K��Ѽ�@b�-@�	 ͽg���^��2�S �V-�ӳ��Zd�ن���X�>Q4,f�)"�)�ז�]��� z7��V3Fm���D�-�b�Ag{F��L�X,�ݛ�sӯ9� �H�<6T�`�n6&�X����Tw�K=��Sl�&� �E9�hc#���r{�_��INkiH_��\�ލ�c�d VY-�����܂ɞOC�TH8u-�S�[�j2tp�|{?p�ą	����t�u�6�G�,�� L��[��h��w#M(H#�𣌕��1��nȆMV����|�6�C�Ł?�H�%X��̟P�F�3~okx����\3:'ec�(%%%)++
��Z��W��¶�xdT�R�����R;c�K'.=�Rz�6L�o�M�A���W�ñ�<��A[�=n�;��Аz����=>n������D��a�T�+���(�xhQ:<�O���=W0����������Շ+��`b�.��گ��2����_b�_�}�:�.1�t�@b9-w�ά8TY-�0�}�*��}�Q�w.������$!�� ��	L�]���-wqFD�DyR%`V�z�un�~�TUMZJ�oW�f�6*l"�&��H��G�&��m��>�G��2"��ډ`%q(ͭ�q�g<�X�6�M_J��ճ���1�{2@�kW�Rw��$�஗���=�W��{�a��2-KΟm�(v�5}�ع���r:�^{�?��f�ś�Wsz���ߜ�x���Q\���	��j>�f�coB�e��ˮ���[p��u�|�b��?#�Z�w��b ��`u�H~�̝���{�e�/�M�W�֧���H���z^T��3H�L�=�_��v&{�*S�u�3�'ϊ__��O9y��h]��{�l|cw�+�P"�L����N���.�����hs���X՘knX���	3z�I�O}���L!�u�7��Z��k�㥆�$�U-5�8�g��%�JS�"�f��;\���N"~�p� 蟒�����s���̕]��Wy�2����]�<T8MR�Qz��z�L�6ͳ+��&U��>���)��l2��n��T�;NL�0�:e�{:�kY38�:!��?y����C� ���<������Ъ�WFh]�SKw"Ub�c��mn?�;$������l��?ͻ�*ˌ���<NR�{�c��I&�u;Ȍ�	~^�[_�1��98#���v�_»�!WX��H� $L��w��Ŀb;W�ՙ�\j�[G�F�Fnu���_[=��N�5�������v�r����^�و/�Kۮ)`@���rr��K;�i�J|dq'�vXʴ���\�{�l����D��K��>M'#X�PrK��g;^�H���mYnm��$����Ӻ��%��|�q���>x�����A�Y�� %��ayk/ݴ6zKk���LY��Џ���/���SA�Ռ��{��o!�S���S�k��|�S6o�zi �eyv�l�ge��$��u�[��ŷ�n��
�#�~�o�栫Ӧ�����CJ�T=\�$��:&�qm�a�F� hf/� UV��#P�)Ÿw��.�p�r�`s¯�����$�V��GCe� rOGS}�̭��#u��W^-T~�^�ϙ�"�Y�ζ@���j�3ÿ1�[����)m��/B���U"O$��q���j���&Z�����K ��5 b��h��J�p��W�ZE�/#���\8'�U�]T޵B1��"��=T�"��U�@)�jyl���<�uT$��?c�,9�;�Zq,�L_�la.ݤ��I]�\�J٥m��piS����,�-�j�gXY��~���Ã+��
�J��i�mj«��@a+-���$�o"J%�j�;�96F,��$���� �IȻ��Ύ��	BaH��v�$�THŻڐ)`�'�%���ۓP �`4�4��X�\�D����֣ܦ}�{��uD	�V	��.b$��!�/nXrX�-R�]���G+�wC�R���ꔵ�Ea4Wn���P��+YҶ'��T>Tj$�eFIA�Og����LhVK����J��G��d�8��A���u=�#��\<Ϳ�j#5��Иc	��|Bj��M{Ý�?��&k>�^���faa2�J�^���z�Եo�M�f���LlųC
�~���/�l%Be�ĥ���A<X�L�=��ʐ�܌�1��TkM��C��nF1>H����T��ƕ���k+��:�Y�=�N��؈`�n�����!�����v����0��D0��� c5#=����tAj㺁����1�|S���TQ�Ș�|���+Į���gf<	�F��B(�$�
��uE36�׵mF���T�fd��܀ͱ���`�I\�$[?��c�~�I��$�m@�k)1/o�_�OJ-�,jTu��ֽ��&�M�����h>��(FW����8����ʃ8n�7�K���i'����)��n��do���ٻԅ�FS��ٙU���`q���JTF&���V���\�!���N��VH��EE��j��m�Ʃ70?�?I� ����7YD=Pq��=>���P5%����h&y����?M�h�n�ï���6���s4	+�����4�����R�7W��(��B=���*��l#|���5&�F?y��#eS::�{W��qj�3!���o�d�=�U��"_���
q�k�7����4�O�����a�і���n�t-��-�6M�+,���"�,^�"ӍGt��k.��������""D��?���j��?cf�(��t�$͢{�F���C�<YyS�!'�͖��3>����⻤^e��$-`����f#}
 �s��P`ܮw�C���f"Z?�x���t��ڤ�s����:/U��/Z���,�2�@kU�vmc�ƭPñ�76�J��7�1��SH�K#)�x��U�x��	�� �yS���,ȁTϕQ�����m��lO��$�K�c��BR:���ٺ�Ջ=�X�����G�3���	���H\�&��4#"�`�,�M�
֝�Ns޾�8/��!.��������Ew�����y ��<@�>��b���#��������8�VW�νѪ�;q�W����Ð�W����=��^��0w��߲�4��λ��%,�����}Eĕ�Ȇ�	%�p����)?��M�F�:�CD����� Ֆg7vA���P���z|m��'���ϵ)R:��SD�{�b?��a�gR��'���>��wZF���%�a{1�؜�����NވoO���I��9�]��]�T��<}�y(��g0
g�^-v�$�b��C����tD$3�����ǈ�H6��Kh��amJ��3-�z5��GqQ�LS�4��/�*]��k��\�>W���Ő��10��̪����G=����*5x��i�O./�S�u��ܑ�kQ9U���7v6B
�v�xTf5�|�{ ���!��C���
d�$��fPC��r��=�VAI���Ǐ���?�E>�J�]���+q΁�7���۞b�#V�AW[dn�'~�z���/����|�]�3����k�s�9���Wx�|�v�uz{r �����>Sc�1qÅ������ή]a_�yxu��H]�H�9SS��w�/�h�.�_!��@NS�:)���;/��=�/Q�aA֐�m��
�7Ʈ�V{�&��潶EpQ��%�<ÈRdB9�<��b#V�Fol�	�;��(�C����n��� �8�?����x���e�ROFO�g�H�������"q	Vi�HzFFd��L�>�b(
�{�@Y�c!6�ĶƷ-l��q)�ҁ|t�vLٳr2���@k�6⇳�*��	�����V�i�x=O70�p��|�N:z�a�{6�r1T붐aƙ<`�6�Y!���kKK�]��(�a�f��dm���x2W�=�±�i%��o
�'H�-�<���A�%�<%���sp?h�����`A>B��vDm����
,SwҒ�����m��bd�s��{�e�A�V���7ٽ�K������%{���0 3�c�O&
ԃ��w{�{�m�@8�;9P����J�ݒ��$b��f�Ǚ�r�@��_�b=(����� TȜ;$�5�tE�n���X�j�m��{��	��Yu@ߑ���Tm�F�"�)X��d��2�G�m�R�+��(G(+�%R��{vR��Sg��ѽ�T�8�C�f���nZ��jB�[�N*G�棠����8�%|O�܍֋�����m:O�_6�̇�]�r@W�ݣX��e�扲��d^���� zǑU��u��e�O'�gf�� �͏�;e�1�x��+��}��q��%�2*H�n2��J��t��y�����g�׷����<�@�D?V\�p׶�+��%6�L�4�#J�Y^,�v<�_RV��oL���8�]\\�G�e2R���HX��N��(4��^�CÒ�w��s�~�q3�ݨ�4��a�0D���zYI�7a����]n�����˰&-X�<�UpV|lz����*��G׵zh
�=(4���� �,I�g\&���RqA����n��=d���&������s������DO+�~��#��ض7�����3��z�y�Jc�~6�LYfbh�G:`]��G��)���3�-��?K�V~��/p�$���:J�<Z���,~����d��}תC�f�d�帤�H�!�Y n������2�n�$!����O�D��?����W�u�Bp%��fXd��F@>`�Z_7� E��LC7XANC9&��tm$�!�R�iz��[��a�i��j�:E����Mhʙ��s��-�qt���č^ ;l$w���E�w����Ë��߾z���fm�̻�{�e������ە0,�X2�f��cI��s��Z7��[WT0���_-&>��I|�ߡ���~9`�,��,R
F��g�Ko߃�%A���<�E��>�#=O���Uy��͵�Ll|h��oxnwͅJv��b���	���8_�[;p�4����.ɸ.�iA�Y��g�VW����._�2��,���`� չח'��o;�_��P�����b���HFʹ�nZn����R`1�>�G���}/���R:yh�TE\4����
{��%�?���q55T��-�!�>}�?�?`�%5w��*�7�K������(��	�w���i�^yV�����G����w��:>�!���������O�eU��ﷲ!L��Ϝ�罭����g���d�k�~��J�7���� a�rK\ώ�0�,߶Mz���/JVc/W��z���`����X�
ă��A�v�2��ǁÚn- �% �?�O�y��$�V^�B����XqqIhL6$�U�TC�y�<�v�����J�a�*(�+�fl��z��s9d���fg��|�ES�F�/ !U���+�J���[V�8����҅��6-���h|N�^�@pJ��Q�u�P����f@��(�罁@9�F^���k�:p/wæٵw/ ��j�4����^?���hأ�p><F�@v0�tZ4}Y�fM�ʮ�E5�?�q��7:$�p~S*j�����������ǙN�����XӳNeL߬p��2=�8Ӫꞗ:5���(��V�U Vnn�_�e6WeS_��i��rC��G������}\��Is��B<�t�Bw-���#O�	"c��ԑ��;��s%?
B��}_1�5[y��z��J�*r��A��9XB�gӦT����D��:�_v�p��f�a=��Y��`�8��Rc�˲z���̈́�d�5�Aq�n~������ldy�YDS�A�f(����M��DI���f?&N�3�W�;��o��f�����Pe��hU*xx���	gg�������ն����k ��YDn2Ti�б��ߟ!����W�E�.5tVrj%�	^J%��xa�p-{�Ҏ���U?E�4�����>�>�ke/��oՃ���4�m��Cak��e����,ؽ�?6�4��M<-������U�kkV�'BJ4�׬��'\7�'�]�q��O�x�|t�>�<�EO���(Ќ�x��VWy!H�b�9��%���#�iQѤ�fk���X"���?��v�?C���o���t
l�ZUe�˖��2������Gվ�s# f	
�`�]���`F�D����2u�������[���Q��Z��l��b�����G �o?�9������]�"��#I_r"@R2ž���Җ��aѫ�_��w��.�������1T����܍��=6�B�>����Pl��v^��u�k���U`�j��p#�G����0�.��{�]t����ݢ�R�q��)C��A3�x]��[���@0�v�[�mΖ��v�;�ЏZ�{����w?����
�w���x���XY#����N^��B�̸~8"߉���3}I��zo�`�����L�� ,r
�5��n�LLo�z��� ���_݋W�?>G,����yVGoƱ��4R0}�1%(P~uf&Q�����:�U^�7Un�������>�[6nc��T	��oL��H���;�tr�/������{�p�i�W������T���o��[��Dp�L,����l��n'��?DkKze��Go�0ﭭ �<Y��ؕ5�5oo�8�kϾ�-�+�\�)��d���	���́f�p��b�II[;\,��z4�N�_�gP��i]�y��Dg<�	���ho?�+��-��*�#�� �l`Q�6��O�]|�.��, ��p'�oŎ|���8�AOC:�4H�i]��@��BL�|/��yV�I Z�O[�pw�_���8M��'�G�h�0�,|��m]-��-��`�����u{1��I�Wa�`��W%{�ɥ<���r���+)GK/�zO���p��b�Z��:z={���'�Ն��p$<Jb�8�L>�j������[�
<T�٣�e_�e�g5�}�����I
�t)�l��neCj�+�Ii�����-G����K����j��UI-M ���=gƍ'�	t���ϲ[�6�+_�v��Z|�����h�k����M/�x��]�	ӨXg�/ۿs��`�İ=|Ue��N�~�i�w� 7!]]�۳��U];׌�X��r�����J��KRTT�����$�c��?\`�Y�J\[�E�`yioL���'cV��CM��;�6�M�4�!֬n�~k�XF�8C�[^B/��'����<�wF�.��t�冘��`����3>l���m#p<
��C�������NȠ��z��"C�~޳m~�7$��GM�sT��f��ħԻ�?������ǹ=�lM�~��ɯ����fP���>�������g�]T�&�%*E��∄�RX���:�@�M������X[0lR�Q%.->��$�+�����cǦ]�ǲs��h>sW�2y&5cC_�P,61QVML�n�]@T)�,���9�Z������ʎ۱��C3Ug����T�a��`D��4."���Ļ/{���#l��ޓ�px�#8�cC�L���A~@��3Q��(g9�::4��'�[���������&Mv�kW��m�=E���G�E�Ek�Qa�i���cG3� ��=՟���u���

**X���@�����5��WZ�A����\�>��\���#7Og�z��Ҟ����A��ͫ�Pw�!Ѓɚ��b! �S�O����c�0��68�y����3��ي��|��b��(�\(����B�+שP��G�x`٠l��������)������7�g}�1S��,���Up��/��i�V�<-�rW`��Õ5�~N�]��7��_!vLL������g���xV�G�hL%)���y�����+'�玻�@r)�"RP�`�ܻX4�j�S����y��%�:��{7w��Tl��c�Z9T��R����h�q2����6�:�j]����-ƶ�Ɠf.Y��r�Ny�O'Ĭ�=�D����*���S�UPݠ�t �8���E�JN�`�2= �S�IO􍒂�j����ܠ�g-���dX���tu�x]@[s�������>���\C���j)�o���H��A ��d0W~�����d$F�+���q��b2��?%^��90��R0	�s���ܷ2��>Vv�����k����M����89���b�"0��c�ҭ�h�k���Z�Pf�&��1�U1g��~��9,~� H�Q�X�&�l�ƭݗ��uL[~�s#���_8QG*��?�s)�ɜ�����lw�6M�V�9ˋ�lZ"N ��R3�m� 1�8/��'�_]'<��t�zϭ_|�)m����4vQ���l�w*���[zȩ�����l��o����O��7�N�*zo���J���]ݏ�������h� m���GD��wv?^�1���o]�osm�>y��M +�:5��}	�������n���?W Ҍ�9@�B��}�Y���E�eC�Z6��-��&�ӂz;���9�Rg`~eB5a5K	���ʝH�=��`�i�9��T�N[��9{�7�)���b��P���#6��?v�_(�e�n+(�V`m7`��]hm��vHݿ�O�fL���gf��� 2��X1_�����{�q���ֿщ��{�7n5\!0	{���".2l�R$/V���wDe|||��{`�e��z@\x����6kԔ���1��m{�m�d>�rr�bq��b���B��9Sz��(bk3A�NM�d-��U��n�	��;�����Qx ��F"J2���}uOY���$�kwE�볉_N[��G �a>�@��
�B���m��6n��i`�����t�t�o��="�᠘	�ֵh��
���p9RX�Fr�����MY�*O=0�L�wBT�v׍����QY�4cF��U��X�� 9xU}ǆ��(�����)�����ɷ�zv02�"̩���v��Ӂ�b����x�	P��[��k�w�ݰ�݅�D(�2���IeRJVLa�{�j5��Y}�}�2`�%� ����U�|r��f�K� ��g(���s���@=§�a�Mg��5~aɛ����e��f��4�F��愊+yBU������+U/��咵L&�9��v�A�ۚ-�cY�g� 2���E�@�=)�Ĩ7��j�466�?D?��'�elȄ���=�&pŒ/F]$"�X��+sa
&ކ@,%���<}sx��um�XW�nW�]mo���Zmc�����նV�z�=���W�&���ƹ�9���8�CU�ף]�~æLۋZ,Ǻ&��"y���.�jPT�5��
�ɂ�K{h��A>�ڴ^���V�=愂FZ������nloדs����h{/Z��9�.�D�M�E-���#�	Gr��4;5��Ӻ�>WXpI�J�ڧ7i�����]� ��V`�D��]^O�I�>YWy#X�.J$�K��j��H<S������r66����g@kK���!%?��4�
���z�K�d��&t�Ĉ9���Іꭟx@?�ى�wU8��;Ĕ�y�y8���������? ˞����幅QǍ�#������~��>�&U?>��uxܰxݟ�<=?�LK�z]t���(O����l�:yDɿY�jR�b�W����z���wxI�,��_��\�t~� �d�B$;�P�Kh��Y��L�׾5��.�K�g�.����v�n{X�/��z��K/K�Sg�^�.�i��|�j�W,��d��aK�\���t��}��<�}[<��'ߝ�jU��o.q�z�����6М�ڪ]�w�@��E�o��t��<���Z���dǗſ�9łꎥw�6�Չ�����}���w�j��ZF���8U���@�ђ۝�+��߱w�I�ga4<�e�c�J�Ik�T��U��a/��
�X��퓉1�J�;�Һ��̰��g��˩�x�)ӕ_���G%��_E�X�bvY|�o	}�!�g�R}�a�E�ě�,D�� �Oo�-��Xvv����=�e��Ѭ����L0X����V) ��a���(������0�ǹ��F���'��Z|��Z�S������:�����s.)i,��n�NB¢���0�����N*���Pd�6�&�^�oߧ�X��t��!�yU��v�n�Fnw� jf0�(���O������5?6�M
s@2���q=V�|~ݺ�,�H�*����gA���Y�p!B%	R�h����e�á����8���G��:��EE����P�'B�Xo��ǺU���%�S�[��GH�U��M������:Y�/�k�ځf8X��<��$�]8E�����!��_R�P+o�5�s�v-����;P)?�Nh������R�[�vc����2� ��j���x$D3�3��b+���.�?>w����;Κ!�绛�ز���O.�mC7y����D&���ޏ��1�֋(��n�����E7�4��l�]���ɩ���8+Mtm�B������=ѽ�>���/�*�<��)�EF����t�c�G�y1���&׫~�Ϋ˟8�M�o�:�H}� 	Ӎ��?��\'<@�Y�����XrR��n6��~J�[M�x���~��`�m���f�It-�]��I����X� �|r�qrfM������ʱr�7���u"���Q�h�L����&27L%��7�<�4��#�NRJ��VY�/Ԥ���O$yI�IF�|0P�	��H8�5@��p�h�� Eߡj�+��ыmh^�jȈ]�bl�=X�js�HE�����ԵX���F~sXh�T3�����	�ƃa���a[�o��D�E
�u �K矃x)�l>���B�֖�����vs�x�Ƀ�*B�^� :�5]����IH� ���q)ڸ8N=�9[ 1���w����J͸�����[Q]�+_�?�	����9�rrb�Nȏ�noo�|����<�S���9A��<��Z���/7�P��(��d�n�����)J��_;�������P��r�+a�y��ne�|��C�+g�d,�t
J��Wb%�?#%��T$)���ם0qf�Mt������Z���\w���ܭ��6Ր��\-ݭ��b�0�l�%�(��w%�;��?��]��H�� Q��+k�AV�r�ӡ��xM���R��~)�{	FCv��2�a{�W�3@��=_�FqC�a�_j�j��y�3q���Ԯ�%�$�����)��i?���n�_"F`��-c=P�J� �N��.�G��>���֚�����9Z`_t/��\�4ŕU���'�g Ua�eXƅ)�a�[�UTT�H��t�lʜ?c}��i�����)�(/��B"P��a`
FyP��7J���oy���/ ��a��u�;8�0_���V��ﺘ�9.�~7j�8�����6�%����bl�R��n>X�$c/p��Lb�](_�w�7�����yVh��Z�g������Fh�l��Mf� J?�����]v�F��K�p���AX/��GP�3��fN���,���7�1�� 	 r-z*@�!��� �rw�k�,�]E%���mۭ~�{���Ϛk{y�u��ʠ� �)��l8��A!G ���󝳇�f��R�c�^F~��I���)ұikX�u�c))�,���,~^�Ƃ#݄�C�+i$�ke�pX�����x�e��(A�`���]���1>���ܮ�("b�b�4�J
��F"X����)�$�����@������X!��Y�Y�[����$ZU=�����EC�����;����6n�����P�;^��6����Pܓ5\�Y�P�'n~b�Y�D�K$�@�����f�S�C��'���m�6���-�H�2z!䱓��;�7]	�����|^T�-f1'�k�B��[���b�j��>ݯ�Sݻ�tK :��� |/�N��H�����'�(ܘ�2�#��V{�v��0��MYϲ�ŢZ�PZ�l����bX�  ��*�MM�8��>m}S8N�g�����ln|� ��g0�4a?��B\s������ؒ��`�������q������e��#Р]�4 �!�G�8�7!���@�x�}�Sҝ2N�8�s��c��6!w_~���X �Ͱ��l/f����Z~A/�<:!�OW.�BO>�(��h��u::����۝&�o�;v����J�oX���]�AVnG��?;X匒�e�`���\ݥ�w�mn�U����+�����$��UD��&���f&]�9F�s�k���I�#�)�����o��H d�&�A�,�Uή}9eÙ�vmS�KI@�rB��R�]�q�7���J��Ks�`�蹂�˽Y�.�V��u/FS���dP���CV�n\�7 ���gK�������������z�,�]�t�I��|�e�5�B^5�M�IX�{ѭ�7�`�|g0�q?�PET�@��~6iI`u���E�I���T.hy$�­��!!3M�c���m�c��-�u� ,���x3βZRt��h�V�)����霹�s��C�&s�����s������P[��>�xޕ��&R+I��%��I�K���J�L���lWo��'Ҟ2{n�d�D��~37�^�}���U��M�X�I*�,?ւ�;�f?����L��Z��tϹE�����6..G�������i78�!�B�L�x���0�=x����HHJ�^2=d1����@��� imR�[�h�0���]�KY5��|�5�9�3�Ps�7�
�x�d��ң�\�������<~��L����M\���HY�#P�ǭ�x��ņ>yx��ha?�/�8�3����Q�^/��)�Gk��1DG�K���L��ƶ�P{���|p���Z6<C�D��1>���^�-���nڍ.~p!�G�2�N0�7�[��NCw`�JK��=ƿ�mK!����������\�<*[ZZ�s�w�>�=�X�Zp<�Z�}�<Z^�\�o�J�#&�L���ᶁ=)�@k����iV�L:��˂�r-�����[���"�/�>>�V�3՜cϊr5�K�D=G`j|��@e��j{z0��6_�0|0���l�0�?�R�UҊ<@�<�o(�<�i��Fed|�l�ۉq���s�A�с�9Sd�z6�����&�+漙)��ݤ-ۻ����/6����1�?4��(W�?���y��?p�G�a��(.
���O//�!�`�;�׾9������ܱw�'�"�x	�' ��~]1�{G�u�Z�s�u��-�5�JE��� Q���N����*�XN�, '�����~�� w��E�ˋ$F��D48�������p	>�8:�,���%~����T�����M����p��_����o Yb�\���Sߵ�T������Љ8�����y4��w�I��6�����f�Q�ڙ!Ҳ���?���Z� ٿ��ŷ�LBIEV�򤸷�{׹B�G�1/�n��R��� b��6.�rF�6�η�'9�P�g�:�y�z��XvS�j��Ag~2ɋ�f�(��+���lݾsl4�\J7V"T���F���z)����'�"���B�A-F�d��]��j�y���z=u�~��N�&�waqx/Q�e�QE'	!�!��NY�'''��RVz F�%M�/���rT��?�M�)8�ڑ!(�v�T2���{�����O��-���5/��|�rخ�Ð'�N,g�_U�(Y3"Ζ���^��\hUTN��W���4*K%��}�\���!�vk\&��b�L����r��O{���;g>��2����ם����?e9�{����c�\������I^��&���/0���A fڐ�����i���y���������-Rm��ؼ��7^����⏰�Es�T��1��+�<Y��iN�)U�&
$��@��b^z셻Y�ӷQ���0��%��Q�Cl�P
�P�r�		߷:�(h9!Q�{:I�Ep���@��� F�Wh�31M��D�0�)���E��5H�c��hbbr���iʅ��4���q���.�
�Z\��ؙ�I��U��J��"�y	���[:y������㾚p� �bnIJª�k�9'vL�`����N�7���<���"h,~��|V����s���.�v�n�R{(��\P��g��k��
c��]�.I�gFHBՀ�[J]6��'��ܡ/m�U �X�y��%G��;&J)�>d-_\'���"0�%����>&��;e��5�A��.	���P'����F�6�
��+e��X}��?����a[�m9��C��Y����j���G��-Nh�T�L��>jIU��K�;^M��p1��k1���vS�����㣅6�s�]^_�~�V��)�Pk��U�]����]�>)H�_�N9�$oAy�W3�9�� -X���N�;��3\pn>�/����Z��I���v��#��fu��w|��1�`ЕSK��@a���
pTC	L���`I?U��i�¶��(sT�����~�j���#=t�S����& ��YT���7�%�m"��M�����ц��	����١?�>i1�sO�t{��2@����������Z&!9�v��BG�������k�(9t<�NHΡ߿jD}rf��E����vxؚ7�^����8��h�*��k`vS?L�/�����_\.tBu�v��־�@�q�W��:�I�P�zzz��X�Ȃ��c�(Ra���{%;�NON�\�*�G���}n��qU�NW��@14��� ����5s��"����A^���y�ؗD��Ӣ���8ȥA�|b��P����_>�?zhzs7QJ�U���������F�eЮ�B%�m_(���Y��G�7x��k�'
��zC*���� z�_Jb"���zߝ���?���K\7 �X��Uϖ��k�d����*���I_R��_�w;�n%D��a���N�Ʋe�+�2���ޑ����U.?��2��F�����-��v���%�����uY�Pc��X��pH���Zgv�c�Z��!�7�_�-S���R�����:a�戥q�v#F��=�`�kZ��\��i����i��f��)O^�9�=��[ߝ,J���6��n@%yV���Kl�����.:�w���ވ�w?@��c�Rg��RI\iM���Ҍ�S�Mĸ�[�H��M�s��,��3bk{"=�w��f��-���y g⊑S�/8����7���@FJJh��ɉ����Tddd_v�AiQkw��=]�=����;��E�-S�ߪ��'���j��/�L�T�k�~���#����Y��ԻDn� x:Q�e�z,B�sE!Q�Z�S��/q�G��Z�	,wOpQ~iE{�XF�l�M��'����5eJ��g��q�������0C��A�4_������p�F9U�jiz�,q�~A���;ބ֝�d���=��^�ф��[��w��&}�e�%�2���+.;Vo�ϲ��0>������p{��n�k�]���Uj���CfN�[�Ǒ�}m���L��ZZx0�� V�&��˵:U�p�ɗ��}�V��A�2�,=����v�4�q�p�aHO��];��l6��\)�D���`�4���H��f�㟔4�G-���@=��O���g�+@� �{�{��ԁU9��J�I%��\+��p���B�?=O�����*�4�dsb�!���/#��V{�E�8v��.�؛&x�V�=���F��RM�w."�Ǉ��E�ZrNת����}��h���{,xb�6�fF�r1J(�Dhtk6�ёܤ#=s� zu'9�- qH��j���M�Lt���Y�C1����/��@��ݏ1㽉d�G��&B./�8�>�'_b<h�T�ǖ���%�N�Ƒ�nv�&�iV���z&�X��o��H�E��m�~Y��-��י@W��C������?Q8�O�������= U8���h��5!�U��s:֢k��"<3��[e[���"z�,��l%��}
��8�Ĵ��}�əM	i�4�k4Z�ߞ,*��\��TJ9H��/�x��Q�^��X�A�k(xq�
*��9,0#}�J�	�㻝9����[H['���J=К�\�68p^݁�a�m�El��im�]uծ��T��kUNr����K�;�Ƽ�{;w�U�t�k�H����4+��9%�=��!!�V���sࢼ�]����p��!��aBk|�Nb(����Q��]��aFE�0Q�Eߖ���w�⣋�}�5on�Z<z�K�V%�1�ZLdp�8��7��IEī�_,؀>�A{�|e�?��qW�i{�x��`e�H8Ƃ�؊@���G���{��� k��<��Z�q�o@";{�L��r�Y�Q"��Q��|؏]-������1��܄�>��]�����~R���f�:��]<�H�]R�!���:���,`d����v�;{�PD�޸�&	�G<�!h	^�dF�ڏ��Jg�0�g���seD�V@ls����Z���n������O���8h"۰#����?s��-}���r���+a�xńb��]����nO���R!���勏��ɏGЁ��!>z��D��ۏ�dz����t�O^D�mx���OVgF��oe[�����#箭�X3�%S���`*�\���.��{SJ���X=�m��T��\_+��%�991d��-x������D��Z/+����d5ٿ�S��n���Մ]�˧���,nx�9z���Y&��E�J'�D�@�F�:=��/���<>Q8ڵ.ۈ�*�U}9YپקrUTrq�j*�D_���u�іԄ�2ҍ#�p��Y��*�4�X����DSOHk��V\�]]$C��9L�vTG�Ѽ)��v����*c�A^@�a֩B�4k���w�����$�O���˟L��H�\o���ܫ��2[�sKZ�e�E����qp�<Շ�H�$%�^�q��������Ɗ��Zr�?���H�|L�/���	��Z������O_?Bd3��78��4Q���d��h��v��e�{�ofV�������ܘCnЬ��)iεEo��Tc,8�!�dHY���SO�'�Y�e�A:@Ve�B�5^멯v� �YL�i(�Q+wq-�b�ߊor�{ɌfX���dldqK�jp~U�;�����Oj�O1���O�������,���D{�a�"Z�#��K�<��X>����E��!!�
T�\�U��ot|�i6�?z�X$�ux�-�Erl�$��Lϰ��!��wžWH��ۈ���o��Z �Y�o���)Ō+H�m�2?+8�A���l���}��b�߷��dtQ�ml"����v�z��~Taq��t��c�8�&Rz�Ԅ����*���sjs[��_6�X�+sy�u8U�vN����/m!a8�.C�T�a�>�F�a�ܼr�Y-����E0�k����&�S��]X�IW�ff������{ݹ�~�/�`�w_?1��&�ڭ��>�:��7�=��_k�?n���(����>\J�T �&8{B��E�.b�1~��'���o���_�?run��%�԰��������������nPi)�e�[3���%��0�_��T��X;c��{���:^�I�|+@��;�tJ�S�؍N�Ρq߈6��"��	�!.S�k(�E��L��I���7��C��?6xZ�/R��5��Q���P�"�9Rm��cS���|�Q G�N�~7H���^ȣI��A:�?��R`F��-�� ���f�V�]$�&|�Z�M�	�`�~�3e�ꠥ�"c��"m��F�a?猡��-:���Ai�c�QL���`;u���7-�W�OHܷL��ߤ���^0m�{��7�@�'lW�|�&l�L����s����u��y�����i��vv�J����P��
�M�?�M��%���D���Eɵ��ح�[�x��7�y�h�'�)Bh��!���ﰕ��X���gY��Ƕ�7���Hx6=/brZ:�n!�B
����K`��;����`���}���/�������lfϬ�)�65�]���'F�Ƕ�Ƒ�l�ԁ�%5�����Q�=t���K�[{����N6��~<�o#���s���{2����Џ�S[''/s�E�ɗ��������Ԥ��C`�n҄|��u�x�[A��?�����v!F?��0�)�Ճ�L��v#�ֆD�D���}�����I}�n��rQ`��؟Qy�xv�h3 �Be_�Z�d���'���;a��[X�eSSb���a��u,n�(Min��x���ؙ�nf�f��u�/�@·��R�S o��'�=�la��s��04������k&vJ4;y	��QqT;jTv	8�����|�]�"8AO����~��f��'3�*���2��	��D_�w�LA6����!���t�P)f�?lx�:���c2���%''w[�1� �8��&��3����'Td	��E�f��ly��V\s�;��,���_).=�{k�D^�O#v�샂�r�OSr��؏G�[v��N���[�a��u�67^��{K̶�)~����=��g�e�S�@��yW	&�T��J����p�~���ԩ̺D�c�����x�K����Sv��x:곦@���G+��������`бt��m��F��G��l��o��H��W���}�Mf���s������o�N��C,'	k�*J��H�>�<�&|&�o_@9c��$>��+�GR؄1,®�O��.�<Q ���A]��]�<��?PL-|i7�����r��A��e,M�`L�1f��$��/b7X;�bq��AWm��S@	� �ԅ6�8�u�W�;߻����v��T�3=�r:�~z[*^E;\�P�ͩ�2�d�(��/���͚���/�μi��e�_T��z/P�EY^C�X1;b,u5�n����*���c�<h��i�7�[[��g���g~~��xi1q�Q�5VRqeYfnG��	(?�-��l��(5@� ��`9.��%�n�)�?P�?�ꔅ ���U֤?^��@��H4ȫF+�wZ�e�����x]*��%��N����۹�6~�I�J�P���>���Q��	V��������F�j� x�M�d�ሸ�׊ܽ�	$G���r��B�_=*��>߱���Og#�����lu6o�\�X�V\�s���@�(��ehv*���0k�ՙ)dHݔ1Md��~���P�޴_�U��$w���B{�^2��d{�(X�~.(�sf�NzbCj�u�=�$R�/�b��� $wa �d|E��%ikF6o(=4^�
K�c^��G,�u����`_<��������A̯M&W��nJ(��1��=��F�)�����Y@��X5�j��ZkuvΚy?ȴ�W$>�� ��X�@	���<�Z��LLM9�#�D�(�>�+!�d�
j_;�Y]��7oX�5t�V�m�6��u��|��۵J� mY~�v�V>��of��	 )?�Zԙ{�5�,�K�ĩm�#g��5lM�A�m�	���ss<��������������FZ����Du;�Hzm��������i)UVBRI��R��h���w��ƫQ� #��V�PԂh*U��(�M�����Ѱ���w`"=��l�������(�R�v#�e4������tQ�)h0��z�̯�&�M��O5�����.�W{n�e�3���?XKŽM���`��UA������TZn����}��P�F���@l����g�Qt L3$�n�CnZ�0S���?��vt�6�ZcE���¼�$[�x��C��Β��)�r_�#���� ��.d4^���{�
�~�>B���Ztӡ�	��G�9�G�^~{��j���B8$�9��A�	�j����vѰ�}��B*T��õ����PX�)�̎��K"1�Z��mA�R��������Q�q���ߙY�Z�&�3��`ہ���V��bޞ�92���#Oi���ڤ{������n�X%8�����53�y��R��JL^<�^��׳�?q�|����tgv��3�/�.@��k�~�fM�x�X�W��$Q�ܐ���;��٬�_ A%@��c���rJ����Y�.;�����^^]�Vj7���V_,�A�6�̓K��:А�Џ�a�����>k@zQ��S�"��kWKI���Ǉ��	-<~%X��_.���F@)�|䣘��x�s�\��ωJYPY���2TL
$�����:4�G��H?���sD��$WדSO�-\�����,���͖<�Τ�q�0�f]��H+��qC�L����q��ܸ��&ά�׾�4T�gS?���)0����jN���iD�!nh?8:���|��+�(�oJ��D�ɹ�|!pG~��g��q�{O��2�J���=(ڴ�a���^7�%�q6����~_�:i��c�f�ަ��~�$"�q��0yr8��[c�rRwU�Hb��4^V ����;�V����������g9F�������M`�<�r�⾷_]7�e�F,�p�� �N\Ĉc�˵�N�qN�Qc a����'@4ɬN4���W�k4�6<������&����2����b9@�ju0�q)�q�2���m����^_������\-�+ �?��K?�zp^����`O�B�N�U����&ڷ��-Rg�w��k�2���w�O8��5z����Cm�ϱ���B 7E[�e��XλX���,�y�H*	�!��	s�q*�LO��k�j���h-*��BT9��{~g]2��ed����v���K�H�����Cߐ�5V�J����D�Oc�P���N��X�Zr��#8�Ā]�������4���@���.pօ�0�R�-��΁=�p������@��_f�xA�f���߰1|�P3�3���)��}U��ZB��>V���_f���Z��>+��z���2� Y�*C���m��}�j5yr���"�?�s�XR^��W�q!������{�mF����KȪ��QArq����4^g*�����&��|���V14l?��� �F�@��y�X!h0ߗ���̆<U[�|����mk�1>�j��3��	�S �y��1F��i7)��o�;!�#�,6�M����ߍ-��B���-���]�X��D&e�9Q	U0m��.�GR�&m\_��,��i�`H���r��`BS
��Lȿ[S1n�e�M�t�D`���b��Ӑ�Nʇ~_��
b�[�1�k��5<�B��hޘ_��^�;����(��v�6J�e�RH��L�R����R����l>��'�g�{��/�8,� ���I�/�Y'"!i8r+�NK|����ٝj?��0�}���ރlP�W�M��xv���\=R�Of��/Z�*\�0��<�>��=I�&2{ϗlM�y�����Ct:�\���5���s�*%��e2(c�w]�H���疣��>b>KA���E����_�ymE���4[�W���/�z�\6xǋ55�@�����|b���
Z��5��H��ƿ̂���&�)�2��}NBw�8�-�L^�2�KxwyG�z�jlA?TlC7��l���qiT;���xZ�7�9�g4�;��S���r���U�^���QkJ;4�:ވKaL����+�� |�^��(t�V3���g�f� D�쒊��!�1T
�u5@bj^lTv���Q��X��KF�@f@I3O$�&挗I����B��m�Fݔ]ϋ���:S)d��X����w�B3�$�y(�^��(@���a=��9J ۧ.^_�^8*,��%$Xg���W�O��l2�����U6|򓓨�~�L��}~#[��F_4ջ�9�T��+-V���yz����@%�t�
6Վ�1D���O����q&�h��A� �]5���QJ�����B���������]�s�e�1�,�3���x1�� ��h�Y���z>�9ly�5��;}�����)K3�n����oi���D�n=�w%���1�G
nX��Xˇv�|���E��3��d@��w�b/����ou �ZPh ��e�6�H����V7�R��s8�qrG\�͖;r,]��B��q�n��,B����c��2�%i�o��:*n���{o޻�rޜ�;Fx����!�{_��c	S�(ccn�(C�ﻲ6R������4{Є_a��{�a��#�������ԶV�{�T�������7����)�4Z�R��~�]mjlrړ^ksEv�L�(���|��طo�bN�X7x��	J}G����<"� QmǙ��f߂�jC!�F�F�wkT	�*������Y:����<��u�"�,����/���ȟ�bĞ�ořɸޚ����-G��6<�%�d�:7���1���^�*~�]|;�0�x��9�8
t��Z݂;�� �N���j�!�8^@�:sw4���� �>ݰ���u:T���S������s~��o]�c�o���=��/M-1�GWߜC��\� ���O&O��"��8Ȩ7���%m��D����{�F���	���H����na�����N��Y\�
O]Τ�p�'�j�u�O��[^����e�Õ|�i���3��.���U�g[�l�P�#@t�m�~��}�e�ub���Dk���Z�������;�6g~��5bp�Y� ܨ���@uR>��DT�Y��@��{�����v°B�#�m�{�P�? �j���ֿB�b-���:���Rl�r	Ņ�T�Ȉ�j��j�`�4�����Uq���<�'5.m<�S���<�B*�h�ls�|y7�T��F-��l�1��S���+/@_?��j9����Y'��-_�2g!併���d��Q��U[�6��l��E�v+�{=�MgP�B G���S[����N��D��m[���3'��j��&܉϶��!��	7�u#�N��-j��
�^�LE�������qG�������]������|�����ͥ4�b��pf���/��%J�q��S������Y�;��&$,���5��&Ix{2^�&q�4��Z�˞���*]# 3�LO�/Z����	�[��.u��(.�Dmb�F{$�v������-In��x/)�yɋv��O�-;��W�����h�����ubb!o��*~��::�V@- G$.q����#5+����Sv�KD��;v$�`N���0�\���.�h	T�|�HE'�U8���)�&*�D/dO�%�MY�	=S́J������(y������u�� �L'�7W&20B�	�rh�sm����ّ��a�@�?�8����|8�~w�Xڳ�&��;
�<��K��C�X	��;��p��c�|mj�&G���mT�7)��g�.W��W�:`:�ErW��ӝ<���g��!D��'am��Mk��Ԟ���t����B�*����7tq�(����Z�~�(�+ܶ�� 9�v�~�ÍA�%���p,*�<
KJV�Q����ٍY�8���e�äZLR-Q!�:��߆F6H�9��9RXx��߿��$��������(<{�����2<S�Vп��pل���$0���9�BѕeP�	v=�	#E-��r�&N��DT�~%��X�K�?*Ƥ�w����wE��rB�a��z.��g�dV���[)썘j�j�Е� J���7�w^� ���2���,ԓ�eEv�L�r(����DJ�&1���ƍ{��ŧC;\h������l��0� M��503Ȱ�윜!iř�Y��X�)��l�nn�;<n�Ϋ�ѩ��v����X �zPPPK�~����yڍ&p����?9��v�^;p�Z���|�7���zߒ��\E6g�7{����K����T��P(߅7섻��3>����/F�x��;W���۫e��@���!2jpʙX�ӥq���\�y9 ��+O����ƚ?�HBK�Z�1>]np^�!"!���I��5��[:PG�ˋ�Z,��??�o�'RXM-�	�g���?��ۢ�xS&,���/?��:o��?lp�`��ܣ��+����� 84SeL�ǵX
9�+��>=����H�e�S��xt��������b�<���.:0����x���>np��K!ӆD�Ժ�;5�W�F�w�'R��OxA�Q���C���R䵸���~��b�	`q�@p�����0�gG��%��xV��,���8є�P��4�-u�@a��FP�vIU�!f�s���������m��h��Q��,26�y%>;�ЩV��v-��A���L����[)===���S���4�0������s��)g�&���j^�T��sK]�J����:)?g�%C���U��p�1Dh�`1���W��~[��:x�q)ew�j}n��ۍŞ�Pc$�W�!��SÙ}^z��1�x���Cr�$ٰR���H�"���0�%>���Ȃè���	$���@$��J �a�Ox8R't�@O/������+�J���#U�=<>p������+���֣H�|D�VS��A��6z�.P��S�*0�it�H�hu67�v5g�����es���_1#����g�[@)����Ô!E����I��
%�@W�ͷ�y�{>��Qjb9��r�?������,n��Q�%��
An����!����}���ik�L�����}9ɵ�9`����zY�=7E]4\�-�|y����E](���I;�Pg8�p����$Z������ Œ��4Z-��J�7�O���`�\��2H�%X?,�øU�)|�t�h6.��R~#�z,�VC	u�w�EYh��E�M�ڼ�R��H&~�� ���iE�m-L=��m_d��T�W�rd�<4���㼮RM!�sE��RIK�_�p��v�7}�/�ʴ���̇�W�?_�Ln����W�[��0�(�C=��:�22�S���߃�����v�c����9�?�y2������|��H%k�8��1
3�%�c��(m�ȂJ�U��J���~�T;��؄ƥ����R��8� ����K���'A���D�S�(9t	�k�uPߒY:�ݘr>e��og���WGI�G�$�fbE�J�q�q�~�=o�7�1�\.ʮS�ճ�¯p�� 'y����E��sZGBIm�*��Ԟ`�X�{���1,���7�W/Ғ��ֽ��&�S������b��O��b&�e���7�65�T��9�ޏ�6�e6"���p�]$Ȳ�	��g{/�(V2�&�͞��6�m��L:�&�;tX���	~=�s%_�<T����Tt�����6oZ�^e�@H+���0ܞJ��Lg~�e=|ټ�.O��0hAK�4����ُ��Wl{���%������Ki�ɰ=�o"��s�����nF�]̃��Շuwgp��|���E&�7�k��Ռ��c��X��f������#嫐�w3e��Ǉ�.���7�~����"4%�P�@\C��h��?��݃i"�~f�
�t��*�l�{��-a��\�3�'��)dT�_���ki����0�R&��tE�s��v�����n�e0�Q�׈1��[ⶁ��?&�&W������u�O�-�������g���_�@��&��l��"D��b9Y	������7`�k-�h̛B6�}�~��B	WKA��D�(�,��j0C����n��l?�os	��x�KT�/L�@|t���]���g*8r�<�8j:X���C�6u�^9ee�����w[뻍���˯�*V�|(C��5{�]|�
�(�Otd�;����?L|�1��^�[��n��Hȼ���9� ݤ�����_"Ƞ��W�r})o���@�i��M4����P 4���o�	R��\���j
�.�(B�Z������V�[U��� <��OZ�eWP_/PR�]gQ�]���wڲv	=�N����N$�P�7c�`Azu�C�fo�����ޔҨv��Ο�^�<��@}9#8���=��;�m�w�*5:uk���q]u��������9�gF-�9��ش�^r��:��yĀ
P��?��1:���:N&Fc�ic4�m�ml۶��Vc�M�ƶm'������f%s�u_��g�C��K�r=ް��O��.!�@��iȪh�M1�����@���}ƌcUb��!���k���D�����,�ʣCEn^Ұ����T��|��[�3��Wt!����|ۍ.�ꋥ�
����dBp��S!E*S�R�.���|M���T4y�����2���U��oxyx��l4���l�tk��S���1ȸCfF�Lq�;���S/*|k�>�O7���l*TD��4�E%�gl׸�暙���q��M�%碇ͯ��CEQY��=��l�gY!'�_kw�3�@��im��z  5�Y��?����z�a�긐TU1aX�Hf���5���b�dA(����@��itA\]�:Ԓ����!�Z��`j��f~�_ae޶�u����=� ^홑�������f������wω��]��L��V��@�Z��z�V^�-�0����h�M��r�Q4� �d82w~X섘�n �nc6���
���ꚩ���V�
�~������(�*��H�	���1s�����P������L��GAӃ�d/Uُ�4�D*���4�/�Nχ�Zj!8E�Tz]F�?��Xb�N�}���H@V���G�\C�'����h��W
x��	��Q�:>b�7�@NY���c���u�C�΋r*c�X�p���0��QI!≵-;�ë8w�(7�;\����|�DǑm{�
��(�-|�t�%%����v�u	:����/���h{xp}�I���"��=R���d��u9���@�����#�
�`�}����:��ȣ���c�+�/�oŻ�NKQ�{�?�8}_c�Yi�Vr�bX}TB�?z�q��WvOA�b�J�)��8q^h���<�w>EW}Zʀ~0�� T{��Sj���/:���ү���en�[�lvfo�����Y�5�ES��X=\�)c��O����g�5L�4�Ը\���?J�t���r��s~�ʼ�Ī��wz��Y+�l`��~c��@��]���n9��g�L��U0l��k"��Z5�l�E�ѓg�f��:�ܢq��A�^�Kc�]�Q�������������Z�*����l�S<�C[��l$f9~@,�L6b�;���g�i<S��I��j���!�H�e�&)�]K�/��
�c��L���d�(�`Gɳ4�ս�s {������������ˋ��#rS�&0�C������J��s��π���J(<�T���^����Q���h���N1��k�	�xi+p�[�֝�_�Ua�:���%���;�C]B���|%/"�e;\����g�����Tm��Op�/�j�c�"��1)�֞I���m�`�3t�;&>�D�-��Mvj�1MF�#��%I;۽B!P�鱎�.l�{��-��?�� �8b9q��`��F]i5	>z��X�3z��~�2pp=}�G\Y:C}�0`5fA|�����q����Y��B��tQ�^�!x�p��pf�E�ݴ����d7Y�K�l1��igT�\>I���[�Lz@0�O��z�*���qaT(���-�} `֪Ui���8r���#�1B�7 ���
��	������f2���*:ђ']-���2O
�Q<���\��]�sF��s�z`~o�o�r5!���9̥�g�����ۢ^�c������[R�Q��?�
{��?<�Ɨ��I�SPP�03���=3�%2�1~L�D��~!� � �/��
���%�oׂ�^A�lд̟K�KsѦ�p�nϳ�	�Q�82�X=.�(��>�K	��J�7p<BZa?�,zq,nG���4<�D��8�8/��2��[g�g���7a�|0ĸ���`�����U��ɪ�SL���}�ne�.��K�v]u��w����s~�SӋ�h���p���x��A<������I���YX_rY$Sk��o-�Hw�{LK��� e+ȅGgp7�����Q�O��(K��6��q�e1৖\���D�����x}�~ха���v�@J�+��d��r�H��R���AE���׭O�x�J�������UL;�%�ӧ��r�=��Ǐu��zi��	�d�m�o�BM��+��)��Qgw'S���m]L�2Ņ���x��6�0�%��	\Q�v �`o����}<��y����A��ú�"��`tevUN��b�7
�9<<�e�=G\E��SN�Rj���m�fo��N���qq� ��t�ܗ�Z��Wy�I�D:��!�����͊&����Mj��v<�ɺ�W6�ykP{� $�s��I��������������55d%������t&��h�uj��׻e�ލ�m��{��y���Ucm�z�-�l����g��}��W��oCȱ��c���jB���ڷ�|��z���_]�6����-X�/Lo�cw�B�'ӣS����p`
Ģ�&��S��%��.SV6��у������[�$���
NlMs�ÑŽ����\2���gg����G�0ҹ�"Li7άo�1�ҋ�l%��k
�8B\�ڙ���38-R��Y:��������ʼ>�h�-���B�J��:8^
�h)S�3C7<��1�z� a7�d�q5Ē�b��/�1i-��a��h|�5�<Q�}2���O �(���g�mTvI���[� �Z�Z�%}$Py��Z�U3c���+"����1EZ��2!1�(52u���s~S�O%e���2s�^�����~Hz�qi��m��;���E�c�����U��f�7�]��k�
�%� �^6%T�s�l5����{�K����nt��ĘYl,�6)Ml���d�_$*�77l����z8�+����v�b�Vף���^��J�8(�����b�w�Q@nZy���>C/FZo�ཤ��������Z�X��*��A�OOu�����j��v����8���j`����;�E�7��Dud|%��H�����Α�yT��-?;{�&�����S�HMCׁ�h ���vG������#�?C���3�7�/x�jx��e%?��p�$D(�_�1�]ä�oy�#�{/�q���s1�DÞO衔������Ǖ��.�.+����q-p@B;��-�-}�Ȳ�\�tkl�W���澹ݵ�	1w��g����޻�]�x�Հ��932�Rs[E�7�<W��&���M3��;j��ugP8�.&���u�K�(!8���{�G5�q
�[8����o�9�c�-5M5U�v��S@��;8_��_������U��3IIIv��L8R��R���3|؉��� ���vMH��9z;��K�a9~��^މ�|�ֻ�Ɓ�!�j��C�����)�(�)�R=�r�mT��d�D-(j����ܗ��n�ӹ�fo��3s�B)����:-~_��I�W�M��eϭW��@�Sw�CF�C�ۓ��ၡ!2f�����=���⧐M�.!�	;�[��L��*�m^��R��N��h�� Ru���o�@]J���:ףj-:
��\֭�E�I;��� #Ӱ����߳�{�:�����t?�y׈�8jE���y}��>i���;��l(7��e�������&:)\kc"�U���@n G+�|/\|b����T�gOm�r4W�9�=l������(l�4=Rw8֡�%l�(�k����{�?v��`r��N�[�">�H�l��F��Q��\yǫ>�`��u!�|�Y�si��&@����Ձ����i5��l���~�㩋���Δ�G�� ��Z����ۿ�[�w}V��`a&���tZ�x��R=T�/!p><�=?t�k���������*���K�N����f�#I�Qj
zl�S�����ᤙi|K�9���I'R~𮽬ŝI};������g8��l.g����4v["��䝡���PXP1�pp����F�S�%�<<ʳZ�m������D\Nb:Ez���0�z+��D�����mQN -�p
��CLM �⻲����J��p~G@E�.��z���ϴR��D[�	��?]��>Q�/^'�s1Ķ�	�J.w�|����[��^�u���4�#ƻ4ȓ�������B����C?Ǧ<~ۊFx��ؾ�R�5�Tk��n�������<^0T:��'N^�a����p.U6c�4#n׬:)��� �l?j�N�<Mܠ��]��޶'H�QW�j���UJ���I5SD�L��?��t/��w+�C�H�OG)GS�^���<H��)|�����X��\�R���m�N�v�W}��C����m���f�$���Bc&��ͬ� ه��ֺ�`�wظ���$]],1+Gc�ܪ l�T�uF �6�w��Ƴ�.���b����"#����&�g��qc�x8��1&�VA��(0��=�h��ּ|��/�?�	�J��Ў/����{9�:���&��Q�X�7���E�s��E��l]��.G�U%�;�1.LQ��O�R���W��$����|/�mK�m��(�4c3�|Թnl)�-�tۦ�����/�*�g,'Êӭm�m/��7 �7����Z��n�L��-��!���w0������/����%!M�H��N��<p���v<X�H��q�yΙ������}&����q(�:RɁw�X�S�}/Y+qE>�ÿ$�'#a�pz��.n>���x<�r�}<�2�xGzU�D�S!��V�!�n�m�� LF��h���řr�@ꡐS���5��P�t��&�/$��������:9�9���?��!�z�yڋ��AGp���2f����؏.�>�o�|��� �aU�x�o����֓�b���u���6�����3���*��Re����r�ړ
��yƇ�Zoǅ#�D��`�+������*�j�Z���]�T��@�1�~2��L��y�.�G�>|O� ��@8������/z�w���Z�w���']�yA�k��3��3�W���4o\��[n���w-�~ s�'<H�q�*�W{��L�	G�w��NQ�(�FeW�Q��.�>��C�ܗ��؇��"�{{{�׻�-v[�L�CQ��]p1��A�mJ�M����FcI_�V��̯�&�0Ep��*!�$�}��v�g;������Ð]�/VόǬ�W�[�����	 $�?�g7����t[�����:�rv8:����ᗋo���H'��x���v[���#�:Г������߫)��'�tlΊf�.�=/^]w�Q��o=xA�r�:���pzn[�*j����E9��
{$1y�������1���~B���`g��[���s�H\-�AHF��v\�I��N��S^[Q-���h�,[��b#A_qO�1T�,�W�^�����Ss�|<64�vA�Jm�ց����Vn����s���9���2cAC���>n���S�G��anj�x�X�>�N����S=f��Jq��3�N�LD�Pcm^q���Tc&m��YȘ!} k67��_��b��z�n$jG�#��8wl-"٘R/�ṻ���:��dy� 睉����Z��%��:P�������a�HT�����O�:�����<s%��c���*���-C�!O�p-�����a�w� ���x��n}^c���N>��ǒP5��/�etK|��ǃre�� �M��Ve�s����<+��G
�F�#]/Q*ct>VYuۉ�V(1
��S�>��J�N:�������8��O��z�ƭ��Ms4��O�\�p�n��؏h���A̚,�u�Zy��Ŷ��Ƹ�xI]�!�:"$!.�рf�>�X���1�'�f��s�i^p4��6dT�Waoj�(<V��bY�)�L)�0���୳�j�V�.o��%ӯ���ѶG��{��0�oܭo�~�لGh�@�
��i�s��-�u;*ن�Y?6y"��hA㺟:���Z���Ӹ_%�B��%掸�~���7`x�,�+��v\�8�����]
���=c���D�֛\i}}�wJ��9{��ok"���9����Ϫɐ���!?��s�U ���[����s|�t(l�K����P��S"��x�����WG�}ڕ�moM;����Ӭ�-1�\bմ�w�ݹ�ͣg:Ϩf��/�.�~�7܋|���g���sz��%C��4D��0ԓg�-ֵ�'���wV���<�O�ŀo�W`��m���^lJ�u�H:T�����F0S��?�͍���0����ѩ����9��r|+wE�u�ޅ}���C�nT;��{	u�2X���༄!}�x5�^d̖{�Jޞ�+jb��6�!��L����<�?���}2��..������ ���*?8|��j2za�����2�O�I�$ed^.�c��>�7�n�`�{�aEF���-�u��*I��Q��U��_��.G�%�I#K���̈́�g�-��{����}{��&���_'�L:����q�d	/���W34�.�(GۊRn���W����ˡ|fGW����{�ߜ8�:����7�q��3Yz�Xi��5FFf�aם��,�MO8�5d����[���&�L8פ\���Iw�������2�"���q:�a)W8%>�Q���=:&O�B��yA�L�N`��*��JR5��&�㑢T��c�$_� ��}�����%w识�٬+�������0��e�|���+״]�[柼� ��-!�O\{F,\��}�vn�?@{���/�؅�X����a��hp��NSCg��������8�\<.==��>��<��BB��;<!���9��@z�-��sB�P�~��K�rҡ@3vYe���g���n��Q�m�ۈ$F�h�IW�n�*��m|߶ª~$3B��" �����SN�0�aéQ��T�>R���1ď�a���,���Bn�T��`l�������F ��ZR�!��w��BMQ,�O"њP����:�������A�/A�B���N�]�5� �P�s�	h�|�Â�?�ҡb����ioTS��Ȏ���`P�߰��;��<����;�;���k���[|<vx�e��-7�;��������ͣ�4��$9��`�\�U\~�k �
9��J��Y�V�8ƈߌ��ݬȳ�S�Q3u���Z��@Q���s����/	xN9 �m����=�!7r���Ѵ'�*}s�I�K�%�_@���Xh��o�h�͵)�s��eڝv�'8�]:j�{swE��l��e6��+e�c��O���	a-�ݛ�dfZ�I�8#�bU���Z�INȠ��A��7^���M,
)��Z���:�@n���U}������f�"�.�7뷺��!�d��@�:�J-�
��_`�JQ�q�h�3�Q|G��/�2a�^�j��t��0�0%�!���ج񀧿� ��tp`M��K5�?[	5�)Vd��`�
���V���V{����(��V�r� �Bt��`��~V�y��A])��q��h�\I������0��,'�WC׼f�������X���[J;<ov��^;��D1�L���� ����u�_�P�i��D�����z�i�	(�5~�������(�BBҌFp2���<�tO�su�ad�b�J��)������9T��:��Y���GlIݱ�����҂U��<l g�ǲ\�B�}9(y�L�R�?qu�B҆�ӓ�U�)����w6$�$1T�Z�:�WoOA�5R�Й���7��5v���mC;b�&���n��U�p4��N���J���t�IkJ�%7��LV&_���lb����K��4��!����K[KE�p`�r=����|�f)>䌖���O�=ך�����q0 ��hG�����[���2�5#˒]��6Q�O�Si��s�����]�jȑ�wU��	�9���B���=�N�s�1�O���y��M��*r彏�@J�ǡ2�o�:�4*r����ˇ<�?�e^�h��cU���9�S��?�H�����m�Xwǝ�~//1?&�[S_l(�>CW�º�P$������}"�v�mn���������|�^L�_t� 뚎k����&��͆�[fx�4 ��.t�8m-}��ߡ���F����7[dЉG
�$%{w�?�RK&��R&�]���I AM�HZ �!���Jm�5xd�n��$��X��w��&E�qN�Ӄs��G"��'�}`~>6>~5�2jg>\i��6��ϴݾ[�WSKq�����ؿ�K<���/�����E�Í���hm��?�,d������U��?\�P��[w ��],:�:ƹ�6W\;�$�㩅d�1�%�<,T��ц����֑4;�r.^w��� �`����|+d􀸙��@��m�;P�4g ����;v�c��/���$�VE�����sDV:صW��	:jX6���2�g�����n|THa�����l���w]@|;W�k����f��.H�f�ʌ�8[#�?_Ȝ����VnsV`A�o�����,P< �Q��c�B|�Ed;��!N��e[ސ��Rk���V0oMK�A�1����}����ߤeA�o�!���@�v|����ホ��T�$�pN��R��3��w}�K����Mύ��@��g*��Ɇ�_l���Qt�>����4��l���P�,��L���H�L�.�#�[r�/��-	
f�@�th�~���&��ה\<f`F�_ג��������t��t�A7y�����G�����u��ұuQ��8�e��]�7�-��Y���]��k��	�j��/L�LHHS}��诤�(@Z��T���Ô"�@ۂ��B�o���oH'B݅
S�#����W��i�OJ����e��M�7��Ŋ�4>o�L�K�(�"��.O��0'E</:C1i�ܘ��	Orcq$����G��U�o�E+��.=j�L�^��/U�0�&��U��*Z�j5&:�*Q��5U���"��=��
�e�g�x��sX���)�,D�(ٺ�T�y���y�\K��n�3��`Q�pl�4�����k�ޥ��Vx��*f�z��!��/�Æ��/>��Ua���g]'Cv���Mˣ=#��H���H��v����pb��[�`�v��2!k�l�-���e�v�Լ�]��PU�"?�tqr:�7��8��t�x[��i���������؊��Ҥ�_�
WϺ�ǅ�����ޣ�]���h�l�>2d5�!�C/�|*���_��A]`6Sm1`N��\�vݟ�F[��N7���_v��I������7�d'���:X�[��
������*.�
I��^��.����G����z�5H�%�Q+�iغG�
��':|M��+fɅ};���yC�fO�?�����ȑ�Y�>�/�x�ƙ�7��
�e�:-��rl8D%9/C;���7�SޙyI�����Y��F���r�mw���KA�������K$�s���Aɔ��j�86�AS�O�s)ȃ�h����,�iKJ�	��4.�+j�^\>��%��F��)�h�:�'��9ܱ���n�܊��Vp.���
���Ū��d;��`���?W�GJ׾���坹���Z��Du!M�� �0l/X�_հ���tla�!C�7Z%�R�y��$���4�o��΁8���^����[���:�0)�+�ӱ��ƚbf�q�5��P��Uk^9\ ��MҕT8�5�B���;9;X?e#���끂�8U�b̮e��:������O�OT��	�J���9�O��;k�,�$獒0|�E�2�c4GF�`��q+?��
"�����nFx��`uV�U�Ç��Zm�L����Y1���4D�@�|ݩ��o���q��fS��,�٫�>�|٧�C�MT?r/8��̛w`�m��t�����P={"A����F&&�4e�W[�%��N��Y����#o���X%Uw�������I��&�(l�"�jӚ�Hǒ�aϕ����Ld���05�O!<P��~}(���k��]���5*��ᾚ�����,X8}8_p�G"]|�vX�|�V�C�W4F3Ո!�N�d�A�����<9���΋��Tzݾ�2���Y/���ް���ۣE��c��������W�|����*J��M���������(kT�M�����S�ϛ��3���J֥=gR�B�Am�7[�e6	�Y~\�c�`���s%���9�nj�[_���)SA+
�^�c�L-�ꈡ��KVV-А�Mr3�3P���נ���G��,93����`���W��ͽ��
�p�'֦�ưkz�;9���D0Iy]l'�?{�s���z31���8w��/a���W�_[��Y��S�����a����pC1�(LP���/Jq�������f0�scE��<���ݒ$<v#�c�IM�1��-�����O��Z^�|O~�S�ܸ@r���+��T���ф�p%�;�3T�.u���;G�!��﫳A+���
���;�'�[:����\�&\T�������.�TsBU�]�w��N/��}�_��54$5�u����z�&P���\.���ԧ��d4p{G� QMMm{/U����su�+ ���U������3����Q�$ik�UP�=Ϫ��p�ԬK�"��i�B�����5��u��M�bbPm���Z��.>w`�nEヺ�@����5FRR�7�R�ombj�	t�a�x|^�,,�j�6�ə���z�����Ð��0g^���cvgk�Q�o[���L���(�9���W�[�Dq���֣7�\ӷGi���ʴၜ���0�W�˅#nA[� ��A�ik�'�����4�n F��v7�Wcw�"�v>�U{{��Z������kJ.oB�8d�fhRS�Ya*?�C���,ǽ�ay�8u�.�*��;�382�B���dժ>/�����D�>)�B"`Z�0y���U���ֳB5Uoj[�`�A�Rܓ���]wS��?���W�[���&�QB_��:eV�.~+7ѳi@���4^@��5f#I��c���u�/���<A��냡M�`�����Ѻ�YG�o���nH�������|-���ҟ�#UDf,�p����ө^P�(xx�Jv�� �L(���.H���^��$2"L�8��T�0]��+mQ�Ѕ¨�h4d�Mj�y����DKM���!�iι��Rt�l����q
���ƕ����1K'�V .>���n[P����&�"P�@>��B��f�w��k�l����j���`�\$���r�� ���Z�g���S!KV���PL6]�24�*Q͍�;�5��|
e��/L\�U�=��u-� O�e �>koy})����$M��jğ 7���`�Ex?8��t�A�~
����Myi�rM�X�^��<T�$#��*�YM�M�K�wx�F��la��a����A�'փI]E(�Y� ��??�RXM� pFw�J�����L�H0���ܧ�Qk���N�X��#���A8�&5�!�h�?��{ra�D$�ʤ���v��qxU�l]w�Ó� <bZ9Ct��p.o��j�N���n$�}:^)����؊�%!�8kw�	�&�����0��s��&nJr������û�H�\P��=Ǎz��؞쳓E&�c�؄�f|�YE%�Z�|<o���'���9k����٘����i/5��P�1�Ú+1�ϣam��wNNN���e���m�s@}g������saBԴV�����O�dxtɺz$�V�tJ �ԧ��t#���/!�F*$ �ZQ#5ð��BCˮ��&Z�P(�bY?�K�Xc�܉���W[Y@��E+Vu*Ҡ_2hhhiL�0\N�
'-�>πH,��/��?��V4�ϊ���v�П�X{9b{EBPbb:�X��~�߁�T�(�h�^w:蓲=��>3��1+��0B-<�D=�L��Mf��w]u�Ҵ��h	��;��(8"}O�ʞ��C?��LS�����hM��RAx+7I6?Tׅ�9��V~��ގe#�^î�P�{QӏlK!Ş=?e�HB���n�p �b�q����{�_zI%��NPt��oh��h�k����Pk ��t�ep���&�"�|�C:,AC��F���Նo.#_�>�췫� �[�ȧ�1��Z
ÿ�=���<���>�~��&Ў9]y���Ep0,iS�BEI)�4�f�D^���͂�����}H�A=ڥ���Aq���0�]*8�y��555�����8:>�����:�OG��	8bu:6��7}UP����)4
V�	�V�7K$�V_�w����;*��-
p�?햒P�A��2�N���E�������b0����vZ�h���^�v�EE����Ͽ ����2�Uh���Q3G�]Һ$�VP7����w,�҈���A��-M؜��ˡ`�;�+�̪6}$b��9��x�8J8C-t�h�է�g��w��'�*B�� K�/�]�o�>���6�=�����T�7T>� �Z��go����y";ɒ�_-�X�q��[�{z�'�ky�4X��&�˺;�.��5�!�0�Vs�a!$�3��^Br4���N�����1�Z_Ө?��*�h��Q�$T��E��D�qA�k�J#������c�Q2jt>/��M�S�q$Ta�x�|��/�����n�!�~�e���?��y�J�:-F�[�
��C"yy89��y�t01�ݻFU�HO��!V��0%��2��P��s�+6|=������+�����|ޗ[�Ġ�E#��WIAq�_��X~L��D�3���=��=���>:ſ�&4r�^���q�\�u@Z����w_v����Dn��8�A��9��JR��7�:�Ԅ����z�oV�|y8�ȮDM"��9,�]M:�^�Ɔ�x�,ܑ���!}��>o�p��1�o��Dny�X���� �D&�;u@��2�"�#7��5�D[K:�]�F�%�6����7�{���T�՘���_r)4��M!�ߞ�I�*��+q"d���?ȍ8�䕉���HO�Z��]��!�T�k�oh����c�l]�	N�����J��`��b�	�״�p,G�osc4�7�ָ�{A���J�ٵ��:*aD�;�L���@�*V1u����Ӟ�q���V_�%�@�DjOʨP=��ﺹTH&oB���|�A����s��WنG��^+�yu8)�gr�oD`��u&�~-��AU�BM�mMJiy_JCy���3����z�:�������J��(�� ���iw2m�z˔K@�8�!xâ""�ٮ����A��oj�Ȋ@9kZ��:������ߜS�<_k�G�cժVxKs $����k����{?��\��?�2��ea}�-��1/�V�N�8��XDʊQ�8J"Y�v�t��J��D.��R�_{'[.�h�� �@��,9��8�ߠ���>�n�,��F�7��UJ��R��ޥs�����u�W��$At��'�Yԩ��+��O�Ң��ɛv=Zz�~6+~y��B|�c���H΍p�j���q|�3�'{�̖���Hv�V��oH���z"� ���g������xX59H5��q!QsÄO`�%�6�F#���B�3�>*g��,�O�*��`�O�
��!��*(97>��!�=7^U�\���3�e��w�J_�����w�>��z#<�����)��R�i���`�P����88Ӿ5��z����50�BX�A=�J]��ʈ=�;W��q��ĳ��il������T�z�	��������&��� h��2R��^���)�HH�y��p��du��mQQ1PՃ"�F1�yD�ȏ;�� s;�Rd�`#�_v���J��J3��^������'���1���zᘾ����^p�_Sy�2u<nGntw�ۃJ�A�_�����L@�Ts{��1�����ק�������q2�os��Sn<xԽ}��\���"�/!f3cb�Y0N�}d�[�A�5�J������i�%�q�Ι�V`u���RvJVx�,p/�H��IG�b_q-۰������,̥z�TEP#���.�n��t������N�X�A�i�z� m`��b|+FA�VJtܯ��(�Va�8�c�/�|ѽ ����X��l\�۶m�
�O�Dl�	���}�pQ;<��gZnI���Ċ���F�E�l����g����"����_��D��79~��y�T�ױ-�<qAm��Jy�7�Jr����ub𿙡��Z���pl��!���K�˃��u�&ڷ�7|����W:A\�1��/�V�	UL�P��u����8j���Q&?�������9F��#+g	[� {R�XA�.�p��-*���Ѹn�uH'�x
e�?����~ކ�����SϚ�&##3�=Y�t����;�C�Jm����{(
W�rŶb.���`�a�����_߅ʰ���V����M�����Bn�^�~�AJ��-}}l2g�w�#�yk�e}3DMtR�'RX�(Q�S��>O/�*�(6�rC��F|DP�%b����@n����������d�)��K!��)Ͱ!����\�W�)H䝼{:�8RDK�d�E��3���|t�Ө}�i�d���`�m'����i=i��@��D�'nY�@BҞ���+�{��o���𳸻kO`���q����_zMW_2�G��8�����o�H����3o�ix�����s�B����5ٟ?��m	�j7!��2A���H��	B댇�?�/>,�\v��@�������*�5\�	��Pq�fE�.���P����q�2��p
���6(Z��"��9p����DZ)��[4<�pE��r��}cHӸ��a��wf-Xs<���k�q�I�TD2<<4=|��P=��h,=@�Љ���Ρx]�5.̫�UTS�݁����\Y\�}��V��u]x�]G�v�����!^)��tK޺�^|���x��K�H�����/�V����H�;]GD ������u�Q�� ��X�n��?��sk�tƭ��^��y4Em���r"���{f�d��=U��u���l����hk3�*gC�~?���r�f�ɺ�1�i�a1@���Q��G�z����غ��0���ƽ�~������*���=�z�Go*Ko��Oa�c˽�d�}D�]ڪ��oy9o�.���_��C�P}�JM t���a�?H�����ф�.8����U��U@��ڬ�P�>���(��q���z@-b�"J����!-���Ԋz�'}�O�rhB^�+M�n��T��C�@ �kE�����f�s>Qc���0Ɩ�InP�_���Sz���h���0��aaJw�?-:�te*�qʫ)�P�0Tx�%�P.�d��j"U+Is2����+�TV>Z�t��2RJ��z�j�y���b��
���pb`7�?����������Y�i+��>CȦdXڡy孋"���*7�qe/�osT����ũP�<y�3���w�C�$,	J��
>��r֏�0�}g�Ұ���K����]]'t5w�� be���B����u�3f�]BAo\��!�I���K�c��F�-b
Q�|#���)}�v]&9��Ɲ����
A�q+y� p����
������Vե�j$Ө��"�`���&&dO?�a�|ߜ���ݿ2���Y���9"~�W̊P��h�}�W]�8���[n��=i{�1�V�\�M(x�a
!���P�C��B4�R����Ys�@H�����]&�4Z����N��Y�����e)6}ШɵCa�|Xx����ۜ+:�Ӗ���?����k���"��lOD�l�bU��M��5z��S"�J��qj��`�/�mn:�U���mEEr�>_����b��T��f�: Y���H�ʾX����LA��+*�ܛ�������x�O�ѝ�>��+�H�l[��G�����&]�;t��쟇�̱cV�[ʍ��e��즺��ݼ:������,Xn����v��	�_</_Ms-`-�� ����:��t֟��d�<&j7�b��?����(�HMj�jo�G��/�Ϡ��.4B���F}��&ga� �0�����p"Q���)�v�����˄�� �uL�m�hs {=���D�L�:I �e��4���C/GO�XY#pb�XM��,^�����"ȋQ�8�#��Ԁ��T�E�T1��.�Zȡ[�GP[�jb������U� �h�2P��t����둌�L�v�\6�s��mg0�v�����1#b �oLP�ωK����O�Z쿺y�Hc�fȐ'�|Z��h%�g�^g���r+�?'�H�}�u���z��H'q�u�p��4jX��!��Ǎ��L�Οa���	S�x��$T� �z'���;�������4y�m�	+��v��;ެ�nh����yf9�ʵ(�rc+�(r!�F&2� y�Z
����yЦ ?@;sV;^���9h'%'g����~b�eYO�������[��W&�	ᑞ� �E�us��8~��d�w��8��q�ӄ��ZrΥ��xs����:�g�Zƍl��s@���Z0%x_~#j�7��,��8%Ꮜ��Y��pב�(P���tPQ��z膡��F�AJ������n������Q������w�k,ל���]��X !ᡫ=��C��F���\�D�ϕ%QBE�����RT}�� �iJ�X�,��y�u}�4i]Ya`�P�,�.�{�<f��(C	B�?�;�.����nlIb0/����a���*�t���+:�����%���������,���ߝ���Ƥ{�v��������|}\bs�B�:��:>	I����������W��_.ǁ�o*D��A���)�龙ڛ��!"�t����G��L��k	�j�0f�Có=+�����fHMOw��?+[�L�L���D53f���7�a�m!�����p5T����y~a��!�-�3�5�7V:ѝ�����nk~���B۩����6��]���K��"2�t#MN�."�(�\o���;�q�w`��mn�%"�g���ӹ�~�ӎ�ڗ��H~���7t���m�^z���$;=�Ec�?m�Pt�6�?a��&��a��'�D0�ň�2�ql��
>� 
�H@��[������\�K���f���b?��D�y��h~�l���	���H�?�p�*�,�yJuto��D�V�.�}�P$y��
m���gz�.PQQyC ��T��(�Ro�Z���f�z��r$�!)]c;����E��Z$eڭ��t�~a�����l��u{�Z�~�Q��}>a�@��=��{�bZ��F?U��&�S�`WaB�d6a��phB\�<����^��9�ܝ���Q�~H��ڌ���#V>Ca@@@��z!��������>��>LݯȐ��.������R�:M�܈����ʫ��C�o@H��W!��d�1nC�al�X���pW�KgH{vM|a$�$�>s�&���ܶ�K���Y���h'�t�� �{"��a���-a�F2Hr;~>�z���%��;ѩ�B�����<f�!�`�h*)N�}i���E_s�ׇ���]E Dnv̳�)�%Ox��}6���0�!���B���w9��I���3�2е^oq[�����Ct��p��k�4� �H%@	Xu���>#S&����ȹYSȞ��$��1!]��^��,/ZH�Odq��=���6�5-�dGq�qQ֦ڶ�.�fڱv�����|�:- 9��/'��yYo�#�\s���| �R\��A5������ǃ�e���	O.�k4�2����{>tPWM:���-�UsſB[����;�����MF*^��7$�������]�?�c�4ZRa�D�q�F�d?W43�FQD�����Nw�[IU�*�-��C�W�d���l>;��B..����)��3��ϓ~�o��h {>?���4e���ԅ)iՏz͂��������˂(�Ӗ�ǝ�h.��!����l����iQ�+Ur��h o��2/)��y�$�s����DU�o�yP�u��(���{�J%,��s=�g�'o���*���bX�ޟ|+���^�B����
)��I�z4k�L�r
]D�����CE�)�Ib�`�6��<1��'r�~�DY��V/�.R��n�ѝ�Lަ6~�c�,W}<��@x�bF���b�۠Z������Ao`�z#��;��=�FV�?�5ol��g���'ZJz�ԅ�`�5�uP��w9rA���QU�f�S[	Ms�N� d�,��Wa�d�S��?�S�j�����>|��H�6���%��#����̚����(ɀ=o�/m:᷌�(;�������'/�=���o��d�_B��6�ssIE�^��6z:&]BBB���}s�d��>�ؒ16�'�X�΅j-�lQ��Z�ә<a�<B�-8�p�n���Gy�q��L� gs�`v���������Q��g�?���7���8N&|�}6j�֯�����#�eI��{�K'�5��)�@�����M����D^]_C�" ���|?�u}��B"�A��'3$��z� M�lۼ/�8=Ou���)X��/�E��H�����S>����n����]�Lr�0dy�X��!��� �i��nW<U8W�q-&��x ��磖nFT��.|c�ye��bG�,t��}'�Tx�dX��J�Kssk�v�J�9CC���沥]��(��&�B������`Iһ䞒o�Ǘ����8V�+�T#=j,�aUmwΚ_���o$��i\����Yb�g̿���z�h3�A�)5��N����6�`�-�e�D\���p��6���I�B�
é�0�+�D�S%�N�b��=�i��j��ф��z/%��Y$�y��ݤ�k���9��$+����܍C�!��P���&+�w,�����*�؜�|]��wj��N�aJ�`��ط{a;�{��C]P���H��p�"�O�m?���BI�L�;0�D���&���(�A�T�KE����xO=j��ꛐ𘕥��0���՟�K�$�)T����~81y���$�m�s�}�hӇfVju��z��Q�F��S��x���2J.��ղG��'9�c����������a�Tl^5 ش����5
o����el��^۶	r�>}?H�A����@�RΡD���^<�@�Eˢ�~��x��\��|�~�_���#�tw�=�����y�	ZP<�W��?������ d�EFi�Y�؛�c�;� �h?�Zz����)�ŷ@S��y:3"̄�5�Z�[gAOL�yJ��xt�7�}��2�f�Xe�Ȫ�<���2y��7�D��Lfh�2��Y����N���(W�':*�ǐ7��Lܷ{C��	�M/���~?��>1��'^�
W�Ĵ1I�r��")n�Q"��n20N��匿�%��x���\���D;[�9ӈQ�0=���Q��)V��=�4'�$p�TW�K�j#٨����|��;t��=�~� �G�;
-f$�Ԗ���=*F��)V��\���"*rOT㽵���Ʒ�J��H��:/{��3C5��'P����x�'�G
��&�GW��f�Y�k�n�s�+��54��w⽯wk�m�n%�T'�]��>�him�;<ߝy?�u������%�rٸX2�ɿ��Ӳ�%xO�vߨ�V�V�����3�o�4s�������	���T�Vy�k[^5G�2�O�r.e�>t�7�~��S�S�����J���g\U���ۜ��4�^ȅ�6�#|x���TR��Ǣ����g�W�յ�c����O���re�����z� ��D��o<��P(0�a�ml�ޘMy�<�TW� ���7@��p�V��{���J���;u����ؑA'�������i�$�o�:' pS���<��SZ�=�-䮏�c���2)�F]���(��������G����<�@^p��|��������9�ؗi�p�U�=��	uC��ly��HV�-��1�RC0�V�Ş����/UΪaL�埪�lȶ�^Q̹nCbj��/l,t�$
�K����������v��!ae�=���w�������/o]����}�܎HD���Ftq�#%l4My�_LO��B�DbG��b+G'��U�Y��C��V�y'S2�gyyY��r�D�Ǔ-�Q��9����$.A$�Ax��̣��;K	�JҮ7�U�#A4�ur��TQ�7�n�\�*���O�h��]��f෵��hJ�t����g�V���17�Q����|�56����6�4��t��$e�t�V��,d?�HF���v��y��F@� ��.��'��s�G�gO�1��\�����q^��A1�o��kV��1M6�k�h�}O�k��^Q��o��i�<V�X��7]���)@J��遬y��l�b��;)g����D��z\{X�'��Bi{:0�-�+=(u�\E��t��#�炂¶m�_�-�����p�_=b~p9w�"�jzi�A�+��9����o�o���p�*/Y�,\�=��`Sg?�?m�p�Ć�֍1��t� w�����"����L>�P$]`r��y�P[��ۋ��}&���*B�s���~
�Uːy��{�z�K/�.KUj��1i{0��U ߂��� �8'�)H,6��C�nl�J�v��=��p�:��n�3h�w�j���� i�vH���3Y���0���ď �?��d��EW'�8à�[��M.�^NT��[�ǩWOaf��C����Z�ӵ�$��X`W�a�h4"&i�S�#"�Yg��=�����K�$ap'\���o@�^Ks��缸v��<B�&�z"z;Y�����v94n��)z�6m����=}��/���^�VR�#�f�BN$X�1�h��_�/f���zH�c�����V�"�=K���*)@Ib11
��ɾjnxD�ݪ���J��F�Ks����-�4��IE�^�S��������%A���������Yf~_�,�N���V�L<[&t�sv���#�)Lg����:�N�)�N8��>��<�������Oȸ�U��	�����k�s{h�T�V����x��l5����D� �h���|�ӰxI��@2��	J0�[+�0��+�Ņ����t��pI��g�޶��$�)�S|C�Oaڵ�8r��5T�]�(O�1��8�
=�(`�A"�f��R�ޟq���r���F�ti#���"�VI���"A�ѽ�m2��6��䤋�H��:$�{{&X�S�)�
E��0���Q��7�ѣ�(�����7��.�v8�!�"�;��L�?��y���{0�W>�m\+�]*:������m��㤐���PPT�n��_n��#4ט�ۆ���(��u_��a'
���/���x��ZF�%�9m��[O��_�~)}�|[�9﬜��.p��)�ߔ J|�D���d/�Я��y�Э����9�pm����#i����s�%�Ǔ)e�;�3;Ƚ~N�U7���n=|��s�mƧv}Jd��1P�lkP��\hϼ��@�����eج]c4�0?��{�*(Q�2M��zx����=���u��6����=JX�2d��r��4��E��QP@��ӆ��)99]&�666.r�$�4�g�*++9�iQ�C�8-�}��?<=a��i׌��!]<$0��K �/N�Ft��m�%�K��u��d�l@�
�+��ŗw�9����jM���݇���+�mc���e��λ�I#v	X��ۥ��h�b$Ah���v5x�3�Z�wB,��*!
�b-?�ό���L�DQy�]$�5�F����~^�O`
��Xsse4�m�:�{?�/��m�ҍ�?ɩ.���xB^�pFΗy�����͜"�׆��F�8�gX��) �R��=�S���f��1|-�b�Y���,y^Zʏ}�����
�1��T����9q���^F�Kɀ����p͏�3k�f��pSC��?�*�8�H�x���Kr4t%H�q2�B)X�9�E}>��f\��˵�N�
�Q��ܙ����M`���M���9]���E>� ��Ų�-�c���{���B�~`A���(Q	}_^[��xe�Pq��V}.���).��$�RRQ}���@��yz��|��D.��/,�d�~� <�Zް]�xL9����qnKw�u}�n����ſZ��#�sMF��N�<�l��_÷�4��PЏp0��-�/Ɣ��G�〘u҅��/h����/͞�h����;	 ������rȯ_��k���R^>(XX��A���Ϙ=�g���q1V
����
�v��P�ɫש������c:A�\<�e{�3ֹ�;q`�Yr����*hmq��tM����1��$��k�������H�L�V������2�_�k��1�Ii��nVD"֑0"XN�OO�?yJ��1Q*�`~y0�/���\��g���e��ֵa:�C�Z���G�W��yl���`��7������Rc�X�1����j*b�gusN+�.�yC����@ϒY�6�c{`*,�h�����{ǲ��ΕV���E����A���{}�O��,͛o� 93tWP�0��[���.	��Ԓ���ئ�ּ?	w&���2I��l
�H��u�i��0����$��-c�_�yS1˶-��9�.�后x�X7u�űqcWEaW  3��yP%�k��?��X:b!	��q�3�5'�ȒA����]n�{���T\\_�\=R�����)~����?r�E_N���;��%�aF���^���+��F���lx	%%,<���0�=���N�!`�D��zmYSֆ�LhXte�&{<l�n�]�	)��M�|������tp�(�D��AN*����^�X��Tv����#�돜��w$�9!a��DCq�P35I��I���1唔>���`R|��jQ�!���ї��hZmmm7?U���P���/q�Z�yW@�h�W�2xU(�Q�K�E�Ӱ��{t׶��ʋ�m��ä́�JЪ4`�4��:љצ�����I�WO��nh2F�3��}�
 �7�B�L�k��1Ԏ
)\nI��uu
�����_M����[ɨ��N�l6�y��"������� �]�Ӓ4���zr�c:�r�#_bY���%*��������(
ȕ,�����װ��,E��fff0]�����*�q_k0��0Fy#�B���|t�m�\�H\��~��#تq��+u���ױ���t�SE�^������iA��cd�ۑ-
�kjR���[���^x�aڎ��U,a��("¡��{����kw�@%ɑ�:)�B]�'���)^8���:��q�h5M%X�	`cc[n�#T��G�о+���3 K��Pg����ίL�fⳋ�F�OL6�[@�'�KQ�s�U�ڳa��$�NHR>�(����U����L�Fv�5k��05 u�qaHX�LL(�����,�J�
e���l���}�3�V�>�S"ވƨ���|�c+0n��K��j��q4���/)����k��qiX�;�5Q2�6aC��z��f�����Y{L�Ͽ]� �*��Bj��f�P�Ï�k���a���@{z��WL'������(��N��;4 ��g�p������s3^��Nv�<16��H�e��]�ɢb-�̈��S�/An��\�5/'����y�m�H�	�����N-���jis�mV.�"M;޶��}�%D�{��zy�w��P}��X6���G`��"�m��n�\#x���=!ݼ�|�.1eM?��f���*å%��B��m����7za�8m��+�G���[��K��9+�H�st�ʋ����(�c���$���fa��}C�^ԛ�kة,�긋����7����{���K|D�
���QG?O�q��m���s n��ڶA7��-�%ln�N%Cb�u��aPf����zv�]�����w�:��B--�p�����"�:��J��0�_nҵZ�pY'�mi�����5�������+MjzZ��DHB)�cJjjРU/����d���r�8���������x��A{s98L�WpF��?�h�[2��#=�����ě`�� J��(�?���aPP��M�H��2`���;�c��}��'	�R@~�]gF?O9$��]��S���g��R�	�-����;��(�!(�H���#��D_g����)���0��n��
 ޴�:p}#��;�1�Vk�*����<�y%�`E%6��������!��I�
�<3��U=+�j^/K�z'w��*$w�x�6�L����=�3,<Js��r�k`<vD�I����@�����L(�� ��+��\�ތ���	8�F��̈w��_Oj:����\dC�"�}�.�?�u�s�G�G��siX�h��_!�F���C�e�,��UiG\�C��������?s��^��ގ���3��{�j3��'���G� ��${��L�i|&AK�l�����&�����~�nUs��^c�T�ק[h����΀T�7��'5C�j/Ѐ��9Y\afc�C?�Zh�C3�w�-�E�ui&_�Q�13(`��c�K��"
Z�"�9�bsn�U��w�UZ=j��R1���X���';y}���φ"�]�:}� �B�����0�vtd�{����Ã��WXX���Z
n
zԘ��Ԭ���f'E�S��L�CC���]�%��9����@�'�B&r�F:�����6���a�_I� �i�"�M��Ő*��+�����Y�ŃM��Wq{���Ƒ�8"A���}�Ʋ�ޮM���'�����2�J��4�XE�9*��d�mA�O���X�n��F���V��Ixy������t����c.��*ͳ%�C��\u)�!�FC~��D�>#�3FaQ��Z\�\��Ͽ\������-�$Y�PS�}�x��X\�mo绹�1��ԥ��ę:���!�g?/uy�	�e�2n�R�d�D�;�s��r#��Jhb��r�t���,�3}l�=��F�������	z~�	�qgZ�0m�jkX�����"�G�cA�7�P#�b���5�?cZ�`�1 �ݾ�N6��0?�i�z��%�<b��\�l����7f@�Wg=ƥ��� �a��ywz����|���z!Vr�Ӆ&�B,�]%==k[�����	��F�Ñ���

��&B �j�g�W�;c�H��;;�����䘥C����:���j��FI�Ā��/]��HKD��$H�*�>�]�L�>��z
�e�k��!3�gץkȗ��Xi�S�}�Ԙ�9<!?����_W� ��*(*Jik,��a������'N� �	EM��$���0��C��fz{�O�Ve���Esy9��ˡT��O��:�T��"���-�uH��9����Vw �$�9���
��2תľ�
�TD����~���,��ЛG�le�E���t������H���й�g��AB��/.�D8ȡշ@�4޲�w�c�x@�d��з|$��Ga���¾�΁��쓟����
>w��ǧ��\�����L��	��Ż�/S-�1^s$Ȅ����P��cy��%�����<ۥ���C<��?`�bP�6��5�UAqQ�Dm�q�&a�^^ݱSܪ��~J��7"�]V�;�����_���|����?2��J1�B�A�yK�P� �#x40p�hW<���k�э��T!�fI���vՖ�x6�e6�ނ��im�	�wj/�L�4x�9o�3���:�Q��%�e�;E�9��4��C �>�xC�k`���AIh�($ s?@��>�>erh�F��X��6#���n���EzL9����B0��OO�+.Hd0TIM�\��Ȗ�h���!ľY���*a��9x/ �u�����>{���WV+�>7Q�Y��dN!_�Bf;|.��}s�̃�#q��ֈ�:��m��i	-�����V��ф�v8�%9!""6ZϒC�o���XI��{Gs�DE6��Q rGO$������R������5Y~ǉ��ݗ�`k;���|��i�c��_����\#�Ϡ�UƷ�pE��Y[�\����p�W��'�y�۫�ܸbd����8��#���OR��'�H:0�ĝ�> �v8�ȟ|��� MKԘz*��N6=��s��h���͐w���#��u���$A��#t���/�w������C�����&�P7Nt���������ސ]�'XxC�~-'��ɳk�e����������Ãt�� cd@��Ei8IRs��m�����>���XjmߛI[�Z��3�r���(�?���f�O`n���S��*<R7�S _�"����_n��PB���*K	֬�� /B�޿�ZBB��J�豜E~�an�=��V*����'�d��u꒩�*��J���L�u��
��z���G��^����q�q��s�ؖ���ϱ��b����9��G֯Y�ML��>�(%� ��|No/lQ�C��m$R��t����>�;$��X�o���>�H	|���ݪ�
�S�&�����KX?��T�P�~b���(�G� k*�Z�İ�Z
qX_�,��h�^~�|d���G�!�S��E�5Bq�@va��ĐJH��So���׷����XZ5�;��,"�"WTT�&��{}�SRS� 񬩭��tf�?˕���@3���^����� k8��>���4J �!<�q!"�q_x{��K��B�Κ�|@�o����I�=�O��N5Q���2ܣw,��M�s7a5=�p�_�f���7��ɂK?�H�d�'+�ٜ�n%Ƃ��t	me��%�2�ЗZ?@B"�%���+�u@q�@[7�,�9�d����k`�E�R]hi�Bl���և���N]�ύ"�}!÷���Vx�Os���$��3$/S��EL�����
����W=1`n����w�dG���s�F م_ƭ�}ղ��w;�ܷ3��=E--��O�p��msڠ�}�����}���'gpS!��J>�;@lu�p7�=l�rn4��U2癌�?���͞"�ɛS�Z��!����ED!�o��������Kޙ�>�߿@Ro t��+ݙ�DQ��z-�:����^��uum��ᆻ<>=��2���>����RQ�;������#!�6��E�
�ۆ�[ժL������Y�"����r��N)�2V.P�l��Ig�U�G���r�`����_��5�͉アdn"�5���d��K�}X#i�ˇ)�|�$@E	luFՖ}ޮc��A+�/�$������䢱P��Z+Y!�3=A������8B8$,�p�2��x� e��ӕ��/��*y����p�����]+� B�W�0��p7�[�H��Y z�@��=��ca��=|:ĭ�$qD[���2?;F�� ?�2�2��r�xK�$Ǔֱ�	p6ڋ  ��k��"�߳��w³O�&��.ka��P������LNC&�}����a���i�F�Q?76^��w��>m�3�W�ϐT0��@�?����D�� _K?�8I�&�6T�,�N��hk���uS���*�7�ڧ���w��g���\H�Sص���~7e<��rys�y+�$ɩ�f!����U�;$W�}�偀h�V������&Ȥ 18����-(�<���N��1oA�fy �u�y��x��`��m
���/�i�U�R$Iz�fM\>"	_�������k��� ]PĢx�$t������D7U64`�݃G�,��� 6� 	I��������f���*�*�P ��:t� T�UV2�	��C${��?��,� �9����؄
½u���OW�ZE��C���~���s.-s.)�v��.�?�)��k�<	���
	ݺ2Q��>�P�w2�m%����pL�t��m8��dB}���^״��)�0^�>���_n�QYe?$c�s^�vt��%���G5An4ZzzI�w���_>���	w8n͗�~��Ub6��HLOǇ�l�h�������+F)���J��U^���G3��$�ݳJE����GH0�sz4
�ԃg�i�۶Eiot�0�,`�K���e2���y���a�,�D�K<�Ν��l_�GN��`Q���X�[�w-�i�|�~ī~M{j*�iCD�Fܽu�G�60�Tv������SGXN�/��t�����m��b��"2�9�EM�����,��r,��O�.R��5jo�e}���Fw+�޾U}_\���DM����ߜ$U�M��,�Lu[g���ౠ��eR ����K��?�H���R9A����.�ttI��apI�ԧ�\��0��f�J��փ3.�Ȑe୎ͣ��B�Z$��P�J?Q�W;�&��L�P�e}��\?����������9�	C���������@*�
8�G��<�Y����}i^k؅���/�����D#�hz�8�@NqW�Gˡ��8$
�.~qzNa5��̉�&ǽ�s��d�

><'���@���M�ی�;���s�f������
:�Q��H<j?Zu����-P�u�rϱ�#���8��Ϳ(9�����;N8�!��A$�L���6�~��7:�IHD�C�4LLL�G@ff��	t*JJ@LLLtRE;����ښ�Å�£YA8���ca�[�d�C���c������(����B��|,�*ǥ�AxH�m�Z�b�թ�|����Za���n4uB��}X�N��<At!A�_�0��ķ���-�O���9�U&.�V�d������ߝI�u��L�om�9��X�j0�Z���y�#�6��O���p���<���i�`��肵�.��ty���s+\�� ��Hћ`�� ��|1��	�]��䨅�I�B��볩b���Xh�D��.�f��:N�j�8����p����q���m6xZ��Iu=;����:���K����!��3R0��w�w0�1-
x�W�D 6�#�u�v�/?���^�����^�B�tKd��[[�s�G�^��|47/�������q�ڗ?��!$#K�o$�����	��1��f�kӀ��`CUF�����߭� �aΥ�E_}m�n���#��J<�A2 ��s�c�SC������P$kπom^��ڶ�'���Wƌr��<F3"BdȮ�2�n>�o�}e�!���ym�$�M����w�&��88d�p�eee-���SC�4��\���[�ŋ�Lw�"��� �;�n��M$��e(ԮAȦ�I�ʷ&!t�v �[�=W�;����fr��!U�SFyI��c�����F�*�3>s#~�v6���oj��冷]�)|½�>\�vy.�{Qhp!G���.N��]���0���v�^L�����`�/![�x��y�1%������=���q�'�p�x��'n���� 2"_36m�b�6a/�Ԫ��z1�irʖ�i[^ܲ#������� �I�ٹKEq� �̐����_XS�w��-7:�mf`y^KD��eW:%D��M����Ws ��Nk�T���	�]A�1��4��`)�?}��&���f�oP!���m��/�Dluuu�i�%4��B��~���E�����	�{�Fbp��XW���dX	h��!���E1����/��"r����fZ^%&�eC�.��M�����z|'_$����{p�Ė���n��D,7����hܹ���;�X�iW�ƀ-��3�C�撳�;p�?k�q�^���D6Kf�����O�z5�V2�C���jq��a Q���� Ձ��	���MN��v۷��XS�}R��R74d����]�E)O�~��6���� quulL2����ٰ��K����1N-Z0�;��4���t��u� J��8�&z�� !����i?/��X�F|=�G@iw�w�mN-͸�b}��&����<o�t��ā\���*���J;�;�@ؓf�]��'`z>k�2꒱�et�Є������ �9<�M�ˇa^��xs���g[��-�wC_��:�>i�%N;�}���xJm1�'��>����� ��Y��S���U|��N<�\�_ rÞ��.��o�ǳ�NAh #x�����Uq��S�r��f�����$D5r���Z`�M��Y"c+�a.E�T�F�;,z���o{���ϟaaHX�G�%���T��Fhy`dd{У��8���8��0�����c������q�����Vҕ���!�{C��5�y����lU�6��?�7Q��l��.�d��\���� ��*�Wg�%���_ )z�#�k�Z�H �Z	�=Q���^
���/����<��,����}I	^��^hΕ@C�j���[Ξ�:(�Ë���=y�E��;w����!����Y�r����_����{CWףizdl,*�o���m��p�G>EC���F?[ʓ��SA�I�׹L``�87����\��""9	��υ��U�W���hRy�|�jV��t�Y�|���-r%�CbE�|�3&T�&]��W�~
BD����޴_��r^`E�JF4"Y#7R�xO=�*^~X�_d3l;�4}e	9���1I�ڿ���������n95�t��fKP&Fx�'N��F������kP��tg�NؖS�X(��oo\�k<�u��~����ӹK����E�b�n� ȝ!%�'J�E,B���١�\��;�QM4i��wm�}-J��"�s{��?A��&�{��,ض�)(HB�"����>JK�,�iT}������Q32J@#|O�Ą���gF$,,<U F��������׫�+h����"5�B${SE7
��g��|�Z��M��|f�U�-���BΞ���'\:��i��A�Q�eH��� �����t���>1��0d�+��)�m>ȱp��_��бˍ}"�A���f"A%	hN�h�	#�v��	���*�(��O��� �y��DhJ��/�����d�ڴ���k�㱱a���:�����A?^!����E������� �Ty|lc%�_�����+L���mΓ��"�~�@}�E F4��i���L�����B�M�U�Ga㙇��&�"��p�NjF�`�7��*;k��e����e}z}(�F1V��p��`���]��K���`����Tf�;*��3n�X)���z�;�Y�����oV�P�U���Ƌ/�E��E���큒�Azx�l�)>�&'�	� ie�M������}�s�:�b,r�QS�6;,������]��?�J��b�
��`�������#�>Ά4�&�k ����8g��x��˨��f�u7)̡[�����P�uz��u�����
��Z��(l�8dx@WW���tDC�v�nHx8�-N���k<����槪T�����u��T__�ZI~�2�Ù���8N�1�9%�_��VQ���S76~?Ǌ����q��>-$�7�u��y�a%��ky��m�`����}����I����M�&~��fd����]o&��օ.��k��;���yV�w��ε2�s�J�y�rk�Cy\��@z�B�ȝ�{���&�z�o'K�@8�Pa��҇�������wh'�c������c>B��������#���J�ˋ;t�l�͛A�+-��>1!������܌c=��$5�"��l��_�PD����A��o�����/�����6U�DB���� ����f�}�es ] �K	$�ih�w���� /i�}�o|ݹ��^�h�QOֻW���2��}�L���n�!�?A��'3�C��J�~I	!֏���{�mm��*�c�U5��g���~r���aIkVi�+�qM�,����K?�]j0߮O�0��7�F��@$=.�Ý~�4�	U�i��E��y���O"oy,�bx�!=�h��G��=A޸�֌��P�L@t���@�ʽ��χ�N�p�fЂ�/�/��q$����j_4^x���a>�H�O���d���ejjXlll�?u5�`&�B�����}0���3������z���r�O��s�)�{�����O�`E����o��K���=�~{��}�#�Od��(5�KF�ާ�g�2x�E�Zy���YM\w�Ҷ�+��E��g�|u	�a&�6����806�]�_倠<և����lL�;9E�AMg�_u;*+F��4�i�^M��W,�Z䡔�VP7�|w&��K����F�G�O��R\R�MF���_`iY��B�b���ӓ�m����������0�RR�
��ggҶ��3��p�
t���d�)�a�� �	D9R�YQ�6J�!���@��D��J��׆}�=���/��OK ����#qk���l��o� ��_g�}�%�W�����Bv�"L\`����TS	?�� ;�Ѕ��o�{�g�Ѓa+�}�y���F�{5�~!�_�ij�,����Ib��=S6p�$���B{\�ftgN��lX#6J�y5��-%��p\�X�4Z��-/60NfSȈ��b��`�� �9����Hgs��ȕ���*Y+�x-Ņ�T=���ڎ3�j�۶0�g��3$�G	�t�[��Pb���g��m���QN5y����Srrb_^^&+xԴMp��7}<TVV��$|}������E9��tu)���!�zI�ʨd����A%�@��������#�>�jhY<�b��\�����N��-i��䓟�4����`"gy���j\�PI�u+���Nj����j�g�O�<�����u4�Q͎�*?��	'��q��5�L3�6^����F�/�����O�4C[<*�O�P���8%{훜�I�oB��$�=�Y��C�
5� /S;���o�z���n����qqR�����0*w�=����B�3g���!9����z�����_������EV�tn9��kƊ\���I*��c�p$��C��F#�)����w�T:UY����z���k�on�Hj�7	�{.��+��ܠ���D���)MNB=U.����.}L���.������ag_�Z�Hͅ���D d��W�ٗ5��E���d;6���5�'��t�������_ob����u����G���s�7�`�b��5H�-Yk=�#� ��a;IB��0�mZ�藧X��B@1N/�zǻӡF��
o�>����"��մq*����\�9�ow��#��l�,J�� lPة�D�.4��'��g>@c?���,��-�;����t�	�"�{wwZ?}x8
$�a%�6��A�/� JZZv&������!�v@�ã�P깽���Z�AYr&J�=)�M�c��$��Щ��TZ\�qo�����G�"�~>�-\������<�e�H�q6l�8s���#߶�4J�^�\���ٿ����Y�T{��*G��-*8�*Xq�Wb��mp18�����3��^����+���h���Cq)ZܽP�Xqwww���Ŋ{p����P �����{�e��a&�I��g���9�9�¾�$��K���Su�i�9��mw�><Z����wcNO����,��!�����9lư`!��u��i�ւ~|VT��LD$��9+�z:lĐ�P
��TVV�nh��.���-�l�W:F�5���Z?'uk�|5��~"(3�_D���hi�©W���ĢND��.	&�WI`u4crj�x�]o�v@/¸)��!+
��ny
-?����5��ó����}v�T��T�fGƒF�4��nW�����X�l4�֯�A��QѼ��;�m��ɦ���T�5��=z2ª�aX�Σ�`Y{l�½4	37�EՐ��w؞�?�K=����p� �j�y� ��������Y��B��[
yjV}l	Y��������h3�*�B	���L�i[ר���s�#;]w�FE��3!2Q�#��WM�����ڏ����h
�<�X�
�����6F�Ʈ�QW�X���EDD �����ӻ_z������BYKU����
���%��������%tL~����k)#5�B]&lk68��̖g'����D�9���V�#��.�N��fzckq���r�~��oA[$D	�/�Օ��ukP���������!�	B?�g,�0�R Yb��{�z@���q�"Hf��f#+�+[H�B�s|���q��������\c �t��;���3������~���E�e�,�LI�kkk{7o%sV��1$!RSSo�i�DL������Hzx�|���w `�@~��D�;�"��0��_S�I�Ss�d���0��)�ǂ�QZZ����f�������M`k��y1��il4�T��}g�Va����J�-*�G��h|��+Grp��������퍹�f��tPH���1��֧�I��ͅQL�g+����c�"�����G��E���U���/��6�@ay���;��Ȱ���7���K�q��-vn�5�4t�#��$�V���j�@��s6+���V[}�2��ƣy��́�|Jf\|e�]��n�n�Х�w�ۢNѰ�c�q�96�-�C�4y$�Z�g�[�]ȘJ�\.��/�Tk��O���?����nwoo��������]�{^�r���9����sZW���w��� ��?CC0��d <�.�H�{"2C��o߀��;�Z����Sn����*�]c/'.ܗf����K�#��Z��4H6��t�zQF�.4�ާ�s"~�X�-�����Kla&���[�� ���}+*^��ʘ���9��L0��ծIZb�L\��fz���@�{ܞ����do�Ϣ���q���7����=�W�"~KYPD�֎I`���a89�����}������D���п�AJ�
 +� ����))�QQ���B�`����������R�l�#~;	���z?>x,G�hO���F��V)��	��M �ۂ��`w뙼���f���ˉ�\��x�ݜ_�]�he���B/+g�фW��>�$�4�vW@����9�5�r��_i��G�w�R�A����[�;�8*��c?�+:�k@'L�?;@�}K�Lca98�75�-��X�Y��4�&����G?{�5
1�Xq���ޭ��ϋ��VՐ���e5'LR�QXB^�lz~g�-O�_��
[1�~c�<��Q jA+��*�����s|lE�|&\�K@��#�Z�0o̍<�[����k�l���L�Q&5"�D�z>t"b����5ڪ��Aw�A�/��|����4�8�9Ò���lF�ipe������Ko	?:���X�-�Y�\_\��)ii��i���@GO1�hZ O��=1������&maA�S�w�������6ؘ�w#�V%�5l��)��N��Y�v� y��DE��}�Hf�I[�ӕ�y<]2�1kÒ��"�_(��"����B�n@P)�9ա�mm������X�y����Z�ryf��l������iy�{ԅ1������6C.�Q�ަ�Qfk1ӝ?9��3��:>臆~;͋�ߡ݃�#0��@�rnM��"��ظL�`��:�g�E[K�33���# Ԙ�HO/��'����=''~\�e%�����D�u�'�W��@��6��α`�t�\����S�}n��de�~w݄�."�P&���VT��/���ܳSa����Ք^!O�|�e�v!X���͂�'�`%65���!�s�rt/kMч�N�������bP{�-���=��S�s���y?W�29U@�j��{YSғ�axDsd��8*�m�;7!-�lhP�3�������{�T8�kC?J<�i-�,��,B��{@ś;nV�@`]#���~M\���@����g���1�E��t�K�$Ⱥ�u{�+m����t0�j�#l�_�UQ3�w�ܨ�:���}�j�_��8� �%j��+uA�҂��z:pyE �(===���>tCj;�w����蟉	i77�啛��Á�Q�����<�j@��70ݿ�_��!(�������r�~�9��Qs>����o��V��=.}e�����|ʸ�~����l"J��K����Ra��D,�dZ�M�[�d�ɯA��w���ĝ����}��+��_Qo��KQ�̤?���X�[ ߜ��_�;|�k�k��U�Ir�»ԑ^��}�]�a���x������{W��|b��h�F�$ad/8��x�
nб��o1GG6YYY%���m��sC�������+��06��s\*X<l��+pJ���ޒ���vӣ�hP����g�9$,��κ��6�p��^'����y#HD����ݍQ3!Wԙ{�o���)����"?��o��-�-޳R������U�e������z>uMiE���C�?m�w
�6���(z�w�9i������w-@df��1���.�q��П��c`AZ�� �`����&ŝ*���{�	�����,z�A���axk&�l������c�$>d��[�lBm��.F1�n����@�/�:��m���^�S����m��L�v�f�wX���w��ac��]������>��N����2�@Pj����2����"��FnF�d��B���! ���p�����a���֔0(7���(������������$�	�-��y*�	��q��	���IF�6�$�ϣ�nf��'�+��_Gg^��f{R�_[��@u�w%p3�v&y��iS�3F��m����3鬖��>�{7��R��KE�c�X(~b��K�ѣ���
�3����68)�|�ٙLNG�mDX���*��@�'�u��`����_�yA�2k+�(�)������������,�{�_*�A�����`B?d��9������N=}�x�i���gnm-���ZIee�Y�������������PU����,䖎x0��/���ƒH�U5���ɫ����:��t���/Tm|�H������A�6�C�	q��w첛�鸐$"�z˚rq���f��;YnGpd�aK	�:��|�|��T��Tۓ4�[��|��/06g�g�x��I]�����+�̚���F��w��R�ښ���:~ϬL�.��I��h���Azȃ�y%���%�u?�!p"��&r��I���� ��G�����0�/���4��O��wё�XH�Gp�X�-�m2;4���[�k���L���`�Ps�á��ʘ�C�H�u:L7�W#7������p)�����(Z�쾡�ݬ�>���C����`�ͻ�����U�V1(g�+��r�FS��(hi!|yy����Ǆ�=Tkk$����0�6����e���GGG@�''��9�g�w�/ �����
g/́�l�8A�!l����|����ka�L����[g5���?3�:�-/��G��Єy��߿үv��j	w*�8�iC5�	�>C0'Ͽ�'?O#�GY��_�����lBj�����-� nO��NJ���8��Ofc����+��p�z�)1��1)P/��O
  W���/�=�.I6ؘ���{h���-X��.


8i�LM���)kkGH}��R���*����9W����^��Ro>>>���U�_��y���՚��İ(�疞��ٔ��%}*8����	a����#�t���R��z9��������3i8�����-*`�G�K����.��"�-7�-uٗ������f�Ami���M�R�B�msǆs�	���u��ǳB.�����TS/g�_�_15�B#zan�+\&t�����5OR�7.�e���1e���8rH����уW�_�r0��J��ф��$���C� m��Ϫ���Fs�g4���>m$.����r{��68X�r��ℰU��@���BB]��$Od����A��:��PC�I�v
m�E��qp�����v���	6U�%%t�x�KK��������;������p�2%��wVwt�Z5\��p��"��҂����������<���U���MI_�����{rrXL�'N�gۻV�vbX9?Mr��<�r��Ha���כ���=�8ιc��w=�f������࿻��<���x�,T���wn*[���[�P+�
|��`#4��D
�PRd|RR,��g�)+�t.Ϳc��]�{[s�Z��9h5.S�z�'��8��l�`��j�w򬂈�hYeĉ���Kط�u��A5���u�vY����uL�x��a��*t�C�!	��Hխ2\6\D*\	 $�@��LV��E�N��7�3[��O���OO⚗Rӟӛ9(�&�k\]�ڤ���_g_e�/����g��8(�G�V�<޼OOޟ���[<�KKK���?j�	��-��V��²~�25�����k�d����*H�ψ��:f�~���Spr”�,U���ھ%��[^���q�<��	���φi3t��˛�:l�'�	��P�6<H��V��)��h"�W���/! �4�Eez�ڟ(�!=^2&�g��i߈�?q޴;C�ߌ��X6`��?⯝�'���sti裩�O��`Ŏ��+)bo���R��,A?�\���o�M�D�?h��P���hm}���bii�Xإ[y�x��X�8G��Ug�m����)dt<�ފ�N^'���\�0��V��9�R�u2�|�:�Wӊ{�<ew35�����ÿX�tGS~�Dp��M�w�o�c'��(C�G
**�*S2�뽿�]SX���H���`AD@Н-��>��@��7C�v�;+���hU�� ��SRB�a_:/�0$����3ɞ4��kǍV��1���=��*Ԭ������EEi//���|]���P�x��`<�����خE�GE���i6�u�Q���Z��]������c�ܠ���)�������W�A׻S����QgxP�v¯/,��F��8W��^a��[���?m#Fn!f*F9��陸:x<ox�r����t6��2.n�W*��?yu�����qv�
]w"��>/��#x���D��d���ң
I�8���,��64@�NQSW7�}7��t��2��=���$�`o8�D-����޺�к�OF�r6��棟Hœ�U+g.g�҃0����.��Ѕρ.K�B)V��J�*\�@TV6�&���fɦ��TTW����jrv��
���38e�<�ډ�vf	<�m�шC
Y�F%ל>j-d���A�/l�h�sDLR~�@牦�F7�v\ׂ4�K�k�
"��F'7�؆��f1�� i^ܱ�b�����=3hы8�������k��h��_3�A�Q�酘��K���SP�i����ws�p)z{R��4�ի���*=�v/�������`} ��ۚ�rj4Ə�h�aH��%7֖��F�b�����|�x#A�k���+ݚH;$c�N*t������Z�p��Y��g���P�lvni�$M%
[���)�R��y|?)��|�OMIyO�XP:�������foo�.���+��w��P��'k|hu��A,���:|��iM�zY����o|Y�L#=�"Sr���r22�S1� �0�����=�Ė08R����O�
;��-ؖ�L�1�uR��
���ͷ���	;����g�o���G���_�6?~�}qW�K�*>4I��
����2��&|z�����cѸ����p�V脌�Ѯ�m��P)Qz�Wq3�y���u��f���t;0m�"<X�t��)2rH:sl��Z� ��郚��)��'WdRt�������S��
�]�|���&P}�:�����x�1���e�����f�w�?��֧�u�7�&���(6�+���nl��e�ph�Gufy��o.�OU�^�I���}*��)��1x�S�A�,u�6nԋ�8��(�T�_i��֠��I�)I�'���5�\Y��L�vy:iA��v�7#���r(����&�󏦏��`Wt���x�z��P(�ݹ�W6���ӂ���-98Š����ds����f
����{Š�Ϥ�b�	������Y�˸>%ac-)�b��Q�߄U#��85��p<��t�slU� ��Ĉ�#��-��ŵ���@��?��jjs&�չ���?�c��W�F�\����~���쬁��!���"�,��ͥ���]��"��ͤ���=���AՅ�B�9�i�}��v�������#��O����"C�1�ruޗq�x���d<�(=��n+'}<?^EN�>J(��+D�X�b��C�@��[Jg���o{ e`�,���&���J������p)񐡢���|����l����<��X:�3dE&�A�U��ڭG8��-5���4}��d�z3�N�=w0�}�xir�K:&JVV���I_�n+@Φ3%##���7?7���3�^P�\�WV������z��&B�RA
��s�hU38W5p�Z���"U������ݹ�qs�.=��w�H�kʴ~~�F������
е� ��PL0��Q�/B�z#�d��]*�M��(�`�ud�c	��Jd��]��g#�qŲ����V����@R�1�Z<��.#8Oj�n<�
�H V+a�o^$��;Z�2�ZnwRR�-��;����#S�Q�y�`��!9[�ln�
f1�p���t����F��K*V�3��^q��۲�Pv�٢|<�D.1htDQ�|�b�uB�77[c�ЬI,m	�L��⢢`��Cly��C,��s{�v1=�(��
���7�T��|��yߴ�l�Y�S�0�1C�~6A O_���x���?�n ؋P�@Ǭ:�XP��{9X�2�0~�gӳH�ʄe�T-�,�Æ��6��i�o�[��@Z�0W�(Z�މd:֪����IrB�o5�b�:( t��Ё����#�Lٶ00k�4�C�ti-����@Hٌ��?;){����>T�_��N�$�)�0�i�jX���utb��?��I��5
Ԓ�R>q�oim�����7�ol�on&P(�X��gB�d:N� � �i�������$ �a�:F�m��TP3lvg}.ȡ����y1!+!�)�s> ���u��Y�z�]�Ԁ 3��5�	5���F���i�|u^�l@�\!�$S���@�
פ/���.�	x~�u[}ٴC��q3lҢP��������5��O�\叚�'�I����ݷx���r��7�c�'��?�|-O���c���>n���+H�艒P�n-��!�G�p���S��_J����J$���@Kk6�W���btt���,�v=����#	<--���i�4���;g0��ĝ������4�]�����Qg��h�a���:���ET�yx�Jԡtz�ͳ�2��u �V��y�z�%�Lqi�A�T;E�	2�A}��~~����>���T`�nha/O��W�p����!���NNlL��>���)m��c���YXX���Bxv6���5���V�͓�?Q��L>��l$����L�镶�e��*��O��JK�	���2��a%��/,�!Քq��TA�Cd�#�P{o����~3�4����D?k�]0��B� 8.?�n��RD�#&`y�t3Ʋ.{��'��`���A���3����:�$���N�u�3���kW��3o�	31o����F{�Ω6RG6܀����&c$�O�'7^�au�l�.-m:���1PJ9�짹�)�?țs�|X;L�O-';{X����>��1�0᎘ĝo�*(���<|�"��I���
�����&�]G�L	ה~���e���\��<�6��I_]�p�r�C�<j�ӄ`�4�g�^����2�#\��DR��NY'k�)W��'B��Zs�$��;:�����������ۋ��%�U� �X��]�!�H/��j ���`8ܲ�$�t��Y�mi�����d���g�
�����������R!~�pq�)M�,#�r�*p�B��t��fP��ة:�.�[��J2�ĸ��~@��'x�
�y)lD`�<I&b7A9x�-��� �r�W�Z _�H���Y�6��u��/s���Y:]�__���������5�u��8�l��]��i$�u����*�j�t�Q��$Or��ȅ	���p��t����*��7����&�b �U��~?|Qt��P<�0�u0G�
Ā� &n��$�=���y�b��������ox>B및��21	��t\]#</�)e�J��V<ې:=c�V���0X�r������J8�F+C��nz�Z�H���x�"sxfS�8�)o�xm�(P��2�I(K���R��e���D��7[��س;h�S�:lQ6��A��%c��T$���_yq#�g�S߀v4��oa0�f�.�^���01����8�l$��㔵K���y���(��<�,0�%�^5�Sac>�N�i���38���yv��xޓ�?ti�<K�*�v���&zO4�-��J;�K�ݷVR�
'���t��d��V�Y��UX�}�ě�U��o[5B�^w�=\�z��6��ld��������ll?&�C�C V�f����ݬ�+��,��y�2t|J�,r��.C4�%O>B�� ����IvMD ��z��`GE�< �n�/P͗,����.��^�1dM�5R�z>;��C�\���U��Y)qn��UY0�F����*$����7$f4���G+��}
��X��c����,�gG�,�8��C��A%z�Y?�$1!X%F7t�v b1b�qb�b�ab�٧`��!\J�B�U��p�"�S=�[� 1�9u2v�t��������k�����)��5k��8�#p�:U�7w�A���zT��@$g�Z3.�D~�3�������R�,ƅk(������yR�3]���NȪ�ߎ�f�x?B�-�6�`;Af�^�m���UP�uO���<��g�b�3�b>����`$��$dz�Y��6+Bߡ�8!�u��h��a�5�_Vv��f���l��V�J@��%�}o����t꿇-��B+
��N��6���D� ݗ�T%v8���̏ �9�1<7�hΜM�EE�	��|-:�uDdp��e��%���yԖk����H#�P����upZS���\}�Z�hN.�E��k���h$��.m�kk�2+�b�_�z��; ��܎�~k{xÔ_���T	��$��gp~��w�=�^葋��N|�̃4�y/]���q������N��M��N�E0����J����A��9��9JH� �8tH��s��?P�P%B?���}!A-FG�I
�����
��vԕ`Y�y{~Z��ݤ�����؈y
Aؿ�[ᦏ��b�.�sC�8�FɁ���z�����>����C��7��Wf:�8 �!�oo@خ(���9A��"�e�P�&�ݮ�1�H���֢
ƹk@p��5ϑ%[x���ß-�> ���s�$�Fx���6~��v'�Y��r��D|g�rc�d<�[Z�%33l/kB�O�:X�~ ���]��,.B�xd��X��Խ��^����run��H��_���rsH0g�����U	�~n���s�/K|�q����q�;�p���C{�hO����*�'�P��T?�r��4�BP�^)"���S=_�^#�:,�P� (��4��w�k�qϔ�@N:�O�����m��"���HZ�y��kG�GS�v��gFl^8O҅��1 zkB��__Uv�5J*3��%�6�]򈞉�cb�Uh����\�#�hD��y���=
���Z'�w������|�n��C�t�u@e`W,�Z��=��I�_�zik!�5浮��ƭ��Ds�K����J�gdBZڻ�i�_�T-�i�e��7����B�0�]�a!���$��2�?��#Tu��v���}=.�P~c�Ȗ��^�B���K�`j��%V���5Xu�I,�Պ����lw����bU
��Ԣ�4��/
�=�Gɬ�2���N�XAc��N��@tPѺ���ҏC�Q�V�'�6��)&
��p����r)鐺V����l$��T�Z�ɐ� ���\e ��A�����y.o�
���E6��Ŀ�iTM$�+����'	�
�T�X�|��=J���"A珪"�r@ԋ����F����/Vm;,����	J�7�?jQ���7a�Î@�G�Jx�!�#�y��&�
̊������s����l,m~�'x]�UzY�0�%^��_SL�+�?��<�>O q�-]�=��М�:��Ǫ�Tc��5?�����A��Ѿ�6�!~�7p.����9�y�Vg�_�!���b/~Irf[F�Q�����u���+4���3��K�m�2^`!�vc���I�N'�	������?�_���E?sH��>s���D�haC���bd�W�� �������؈8����OFs�Qs0�o+,_I5/�3���{���l<Y@�R2V=�?R���e�+b��-�f���8r�\"4�h���^��-�0;� ���h�i�!�	C�>�α�C!v��R	�~��T.E06U��h�_��zRp�.� �uܭ�������]��)i�,�jür4ګ�]1!*[�O�ŃA�p'|����E�+�ghN���2|as���`�A�a���F�$�L+�G`����:�>��H�W7�o�Xju��G�� X�p��q���O��������|���v]@Vl����|Ou�����4'(���O j<Y�'����F�i^�w�Ӹ� LɅ�"u���AB�U_�Xv_�q��0����6� l�i/+݊���b�q벨�<\�C�t;.S�����f��?���(���K|�$	��MGz/T���+�d�$�<��wZ".��ؒH���~��L�N6Cd��N�6:��  �z)����m���d`���J�Mʢ2��y�8�����W���L��H�oB0r��vr=�>/���z��t���Jpdf۷�50ǳ:]p�h&�8��5�1L�3␥mi�8x��E
��q��5)����I�tω1� �$�]���?8E�A`{��J��mepk����+�K&�K��k���\H����[��}C�D�_p��ii�[�Ƹ�O��뽷I�����۴�1�g�EbC�~�:���Y�\����[�Л�1��3����mB0���	&���ن��E	�1Y��V��#e��ѵ�l�������+��S�V�9	C��i�s���u�(�/2�<yA�*=��A�v2���uAQ���̈�}���U����NY�/���Y$;�����i�}�압���ޔ�1}�~5b���ۀ��d��d*��ۚ��6�H�D�S���z���9wL����r}�(��]�^�2Q�������F�!:�V���"Z�+����j����]��?)�`z��"�yܸӡ�n�[C��E�������D��i�_�Ʈ���1.�G��JF�wU���w_(k���>����%Ѩ6��P��u���\K�AqK�����a��{䒖���&0QM6ȼ�B΃�Ѷ#�*	Z�Ȥ��T�=��9�7v&���G��|'C7�� ���d���b��` �X�PM����(භ�*�� �;)�BHM�%��(A	��}�S���ڎb���A�p�@��_J��{XPZd�-�d�{����`��~~�JK��-��4���-p�P�,�|w5��F�A�A�!N�ګ�����#�9�Vq�{��&���C�F�v��5FM'B�R;:�z�n� f�e�7��'.�-��c2�m�8�2���F�_v 
*�	<�%gT���Hr����G�[)JT.�MFn�\�A�� :�E�Z��NO�����CXT�YnPQ_�����k{
�2П����j!�: ��F�dc��՜?�F�!��G������$�,�~�C!{�W8�!J�<"�:'{"����r@�i���/�}!21�������.i�֟�&�y7���������K_�։�י�Z���ը?-,aby]��w��k�h`�X����*I�mK��e��T���8��Q��&Na�����"[I�N��Z깩��b��f�B<ڃŷa�	��$
b^#�)m�;$�� �e�p�W���ڂ�P9��	�8�,P_��;�a�������q�)ЛWn��=���q�R�s��U眲#��`MET�n��R\A70�/�E�*?r���H\VيȄ�����dA�&u�c5C��qd�[�]�)��)��Z�a�[��s߭G�]^��X��n֡i�g��?��������&���k�8��~/�6��J����#K�m[�R�*��jJ�:���9+��\����ۨ!���iŝG�J�R�ǬC��}Tzya�{�>����k���y���iG[~����)ܾ% ����J����i�n��^��=����S�4�6iYf7���d~o������~R��Ŷs
�tQ�|MTn�����h=�x<����.��)��/��%�z!����ۉ��돰�Ȅ`�z��و�˓p4��J\��
`"E��B𿱤p�[��m��2z��z���N:6���6�"C�}��:c����A���pO���*��0����D�Z.:�}p�q�Z����z�엟f�#�O����V&NN�r����$�o>��,wkpU�5b��39R^^-6;��E96�뀎����rRP�$�������� �=8μf(�Z�+F�$�bs�)xL�Uf�+3�'�ֳ7�Y��.R��q����N���L+�z�;���qU�~�����*?�3�ImN�ɲ���Кz3~�j%V��u �����Lx��x�t�.��r�Ai�)~?�Y������/�)ډ��1.,uM)C%X�xSM�%��?Z����6���o�6�6fn=�Xe��)xke�r��ͤ��9즌�ki���:`W�a ˪%�h��X�7�!�_)�]���`�ú�����k"b3�,����D3݉~/��AO�Q!��+y#B��#�f�;p=E{=C��qf��1ԖrX�[�4?k���>�XȬB���j!�Kp�뭍Ó?h�>?�����YĿ�$k6�q#��}���1����O�j��/�9�H�
������`%���L�	�!h}��E<=]!���1)����&k0�������j
Y�m>��z�y�
Q�o1�N��7oa�O��KH4�M��S�s��kO-�tE�/�z�N%$7Y#�!��яq�Y���Һ���ɚ�+�<���N�� �9>l�	Sjm���^��H5B�'v���	
�#�o�:]��t#���s]O��i�w*Ո5�?��G�#F�6���������ڈJ�#%,=�y?�U�]���Q���Ih��(Z��5O&D*�����; ¾ۇ#)'VW��4^mq[9�H�6��I��u���.����i�>b;��8u���j�#�(pvѼ�@q�����]��7fPѸ��xIp�ޫƻ��Tg�#O~Q�tu�A��w���i@���rzk"e��x�%Y�_	����ʒ�@�;#��&[tG��=���ct��U�s2��Uߑ�1���ɺ��������$e�I.�>�t�N� V��+Bu��a=��+�T�Q���/�����t�o��g�P�6�yl��N�<�{�qhW�	��/<!T0�}�u��o��?َK��w�/r��`k>�V��({}/7����6 #�ߺ[�Ẻ���x�����B}�њ���h5�
b�eG���#��j:�J����nx��76��a��U��fq��A2�4��֢X�%oE=qآG _Ä�ȶ�R�B��Љ�D����k�x�Z�)Ԫz��w�tv�llL�*�A�`���lĩ+���>󌤷�-nkka��8FC�|k����Z���ml˅����������ڐ��.6v�'���(̿�V�����r�����kr���|,�����O��Dޔ��.%Y�ڈ�?#����g��-�EFI�%�w�F��A���y8K���t
�Y�M.:� �,Ѓ��C�L��[S�d���+@�����N�s���WS2o}]'w�N��P2_���m��;�Jpf��xCs)�M��͓����KY�jW����e���h/]� n#�� ߷^w��G �Y��-yg�pQ·���_�7Y�m�Z��UA7����D3)��f=o����d��I�Q�>tH�ӝ޶��t�>���*9jQH��r���~�'-CQ�vP~��[����p��ka�W��v ��5��3y��;�QPY���drU]��!c��+����������8���S��Q�Ѫp^IdLf����nM��v��������)����ӟ� ��:��������x ����I�¯�������%�֋[�i���8�$)���!+��e4�X�W���a�U���I"���S��Y����K��(ފ���0�&j�A��HBOW�� �@��.A葠1:8�6�)V���8:>H��bp�����mǹK���/A�$�o%a4�q�c�+�M���,�&P[��O�e�Pc�ՒP}/-ow	�O-#r��Ǎ�e����KKɋї��#?Ѿ�y�L�J@!��j	A�L�Q�ן��6|�C�1��&'9o12�kX22b����� �p�;Xu�c�Gf� �8]5����l��bH����n��D�%:5,W!�b�~ 4���0��3��"�A�� h��Q�Ɠ����J'�����N^���'��H%nvlP���:���\��ڏ�CTg��	� ��|�$�?��q��f��Éܻ��aף������U�vU�TD�`O�l<8��v�Εbړ�&��|)���E�2�Y���hǐ�����1]�bD�n-V�<�*hr���E]��S�ς�	!��o#�E��u|.�6^(��G�>^�����p�?9}�U������ ��a"&J�C݄0�r���Nh�g���6.�����ߝ%g���q����ɱ�=��6>�Uv����)rF�h�:B�XH�,D�+!5\����B��օ�������-����e/H�s-O�p�C|�.��7����f����P��W5?�k3F�WX���gO�@�db�}�O#�N2�e}��ޯ
�f=�px%)OH�H��u��!�w�w� ��;��ݟ���|Hlk�J'�|u6�-��^�����P�#<`BC�W�:��ϳ���#0�x�q�.�M'A�,�]P9m���_�y�b����B}+��6�742�O3�Z��Ni�������L�����X���D���E����O"V���Z��/��{��6����{�:��AyOb�-&����2U�;�\>|�c�ʧ?���l%��4ֱ�#=Ϣ�c��k�A�=�K�.��YR;��2���ǉ�z�d�@o�2�,�����L�D�W�A�y��ք�d֨i�"$�ڊ:4�ĥ�]2H-��
�eu�����E��ݺ��'=p�����>����$o�T�ERr�*	H�2�U�o����̔�����VT�jO�?����Y��])��p�����D{KN5~��{e,4�o���]J�a>*�Qyk���wt��j���f��N�tJ���n�@�t��/㟉�<&Z�%��bm�!KܥR�TW�g��j�:�n3���+�S_��c�YqA�!����ѻw]+�H��C�U���3Y�1��^@��fW��E���Λ�:�k��	����ǒ����q�B��:�k�K��s(�'��)���UK��q^��<tm��}!�t�75�Ww���fd�ya4�/��4�x:z7)��V�-p��;ᶕ������?�fa��CH���2�r�z,�0b'�L|�6d�2 r�_ۦ����ν�ٶ	X�2��{�H �ϴ��;u�D' ~���j��5$
[8�qK�3fLb55�&���i��/�``�w���
�O>�п��TJG7��7�*��/����8���T��V��\��f�����ԙ�Lc%~��Xe�����&�u�O���Kn�9r�����L����S�����-��ښ�a ��	����������!�����w���>��թ��sf��^�V��Y8�$<c�R�V��\|�����;��Ư;5���Q��Dމ�����.��0�)5��m�@�����l���3^�Aw����skz�j���O_�lC��爭$�0�d.ͮ6�G7��{��xt#�d�x�Q��q����[�W�� %n�i�~)��|�ڨ�<���5�|ގ$d��^���P;�y~����{���"�}�)m��WZ�qи����y���e��oYO�4�J�z8o���0�C2w+K��8��;ɸ��Va!m��H짥%2�L�u�� &
��I:�=���y�Y� O�߬��`4ʽ��
��dɡ�Sv�͍�ؖH�_����(.nBQ�vH����=�)�� �4Az����[W�����F�o<+�������l��6Ӛ\�r�sf\��;�<XS��Q�*̈́�1��
ر��/�Uw"M���B��?���uֱzD;p:�k���1d�%����{�N%��å$�mJ���\ 5��<)ۨ<8*�S1S�G�2�����'Ŵ�3�l�m �B'E�u=n�� "������1��͓P����sd�����eߑgt	 {�ձΏu����<#�t�	��,��¸N�-����5;��~�����uHT�3�2�|�z��_�X���^$57�J�	vQ��[ѓ*��zq�}^/e���"�s��_��������t�VÏ��5���.ˉ?�������DF>\>�ܹˑ��:s"Y��N4���������Qdzʼ�V�Ks.���f��'��J�{��S�!p����&^㻟Jſ�crd~�V� ���i��z����H4C�����Fı��mp�n:��/�O�UАk�"��ͧ�95�.{"�q�T��*���P��P�\HS�����fI
}rm��']��Y3/�_�ꮰ��L�N��S Mt ��0ϾCA�$$�A>Yw1x]�Fm|~.�����@�{��=>!)��ƲL��$ѢUh`��a�$ή��D����`vqP�.��!_��+x;�jn��E�%!�m�ݭ��e�0F����A*���+��y��I�B��pf٬�(F|{O[5�(�`x���v����`� �-h���F�ߋ��U{C�5�\����m�k�C�����}�m�7�om�"�Z�q��a<�r��Y�:���m��;1�r��� �n r��s�'Тپ��@���K��FSSِG$3�v���*��P��I@��3
���Y�C��F���ti-Lp�I��[��$���5=���s���~�ϵ��(Va,AQ��Db�ݯ��ǋ�$��ˊ���7�1�.:�ܵ3�Ud�ئ�������]ܟ�	���4Uv��\�Ý�7�6�ѥ�/P����a<|����Ϥ�:����s���]�/
�4R~(E�*��U>@�ݸ[��K�[Y�ѐC�b{�-hO�P.�����غh�[R�-I�+�qwфi����vI�T��Խ�iQW��l�o_i�m���q7��=�d�=\b1�����jQ���*L��+�de"��dsr'��[��{L~�u~����{��Y�	9(ҝ����ʿ���k�*V�c�7���Nc@(� ��8��-�
-����R��Z�K:����h�0��b��^S�<�0N�5�M�Nq��2�*��A���p�뵚�g(1o�s�CD*U��'d8�H��h�^� ���2�G��z~}�@h�X������D\f��~%ˀi1k�3g���Ŭ���0:Y��Qf����A���_�KiOp�a�6�DAM���2�cq�`���i��V4P������D���g�-�>l�����.��÷��%n�{��%���5�mx�͎}��T#Rn��.�$&##����=��B�L�����X���6SVX��BT�M$����"J�쵐0�������`�|{gŐ�^�-��@����_^,���D�w��{�%z�a�x�����z]=RP�B=��ｲ+:Q���9�S�*t��+���VD��xL��Y�h���<��(i�J<�	5R�l�
���ݵ��^�_/�n��9��p������==�H������92pm�����|�!�
��>�_<,Dͭ����"C���A4�s��a�Jx���=��d� UO����>����+Z?�<�#+9z�7�&��E0g`܂rfar�<��V�ۤ)��6=��X�q{F���3F:vD]�|P{@ܦ�W�@~�,J���:�L�#O;�w�/�^�m��h����^o���2t͆�P���9���3N��8t/�)6��t�4�;(��r�yl��|��z����m�l��V�|�9�n���]��4&����o�����=���?�ق������R'!�t�U 
Wk]���a�,:>t��py�5.�����5�T����(�f�]����[�k�{1q�@�&�YN�HP��p��'{k�ɒ�m�K7��# ��U�R#D�aF:�$3A�j�es�?��\�P�p�C\:�#�%}���[>Q��<d�D��p��x����*���S�ո���c���dA�Pm��R$�z�L{V��U�k�0z�Sx�} �tS-}���q��~9�O��p�?��pMm�������-{d]��K۬�G�-qD� �KGcy1>I��ҁ�r3=9ͭ���L�)m>MP
��*������A:�ˠ0E�n���c�H��̓�"\E�����Kz~Z|�y�=�$o<6���P��WJ�Wp!�G�O���y�,R�`���
�a�x�ыG;=��{��~<[�����a#@.���ԗ�nt�w%�Cf�1c��w͌Q~*+��Q��"�����O��ǽ!}*���'Pn���X�$��[01Ќ�$�u�,h��PA�o��� _��E�Boi$��EEO2�+p���S���w�
�zD�;�j6ķ�*9��9���T�pp?Lo�d<�sMY�	�{N}s�n)77ôA���-$*�%�	�4C+r���x&T�#J����[��+������l�5r�,��~@U�|�{��,�dŽ���7�@&���-*�0�S}����t�S&H��&P�#��v|�GG��vm�<̥�i5�@"�Q����2�6��K@���W}Q�٭�H�Z�/²Te�ҡ��8�{k����]����&1I1$S��;YYdy����g�\}3���*�g��?�G���,&���k���V]�2| Q�6���:@�oJP�VO���T��ϸy7RV?>�ZU������GNW�ߧ�oۥ����Rd�~�Ut�R�ӟ���ۍ�E�ߣ|
��z�}GXbҸY��F�ʻyy�Af<��Vr�>D>��|����qL�]�'�?�п��H�k�"5.P��-�6Y�4��u��	P��A���Z�xp��h�G>	����*�{�3��ƽ�+F�ŵ���FL?����PA-:XҬ����i��=�bDu��r [RH�r�a�Y���R�0��0��27��<7����N�P��������|N�g�P�44"��sT�i�߆o�J�@��N9��A/�C�u�4f�?e��
�����i�/��Ӆ�2�W��Tѣ(����^Uaú1���2-Ӿ.ɝ�:��g���s�F��0�g5 ��|,�Oo=B���3	 ���(k.H*�z�%�9"N%]�WV�m$Γ2YϦ�YVSUI�O�L_��{�t~K�j�#�4���1�>�����E�P�鰑�dR�b1~T]���,{�"Ѹ/���xr������s��8��$0<�Ii�(��a�~R���r7=�	�I�$N���>��-tס�^6����2
x?�)C�U�a��]+�C:�����ɑ�SV�(�m�����y
����Ӭ���Jθ{0�z��@G)�X�l��p��|�loͤ�F�S��{eƾ|��0ȟ}����/����x�{�8>����=�l�5a��J�& �s������n��Y4��
.,N�?��� |��!�mS�p�����>�%��iv�����0t�ڗ�1��� ?-F�r�\n>� :�r�Q�^�hF-�C�Q��D8>���vS2�fZ��άP�`��7U�p����Žg�����!��^��]��ކ����҇6'�]��	����&��:��6���He��l��H�P��̗����r	�^�;;,�j��]M��;q�E0���M<���?�1q���ɝ�:�Imz���Yܑ*�Z��N�?��y���hF���W%[=��`�q��.j�?��b�I�6�.�)��+3��g��<��^���,\��4"�A_�I����H=�ǌ��U���aa�);��_���ViG�G���K1"�O����9Zy��c�\�S�]�>�mˢ���ڊ���d�?�ᰥ������e�������B�7$� b}V�x�.-��_U�X���O�ݏ��.�x#n-@m�R�v�&��K�W�3uFp��S��bT�K�j&�X�!gh�z�ɇ�ojs�)�!�i��]���C	:xА��bKd��Kr��M�n[q���#N�N�COͣ�Wz�d<�����s��\A�_�kd�rhݽ�ja�:�$^�y�"�L>l�d£����Ε�4�j�(zϗ��+PCK���E+�O��G^�)�9�b�kOm� ����rwߐӆM��x����=�����$lff�9��z3t#p��٦�����,拄
�-�ꙹ�2�l�(j֝>�~^�������\�ȩ�k�,͑�юR�'g�D�[�z��~cb�����?A�J�a ��
Vx븦�����h�5�3�t`�\q%�<͚7��qYcj 67m$F�-��0nP�K5�o@��񈷝�#�	�p�F����*cG嚁fk�?)�o.KC�yu�Q����,�gXPbG��x:l2���.�o���;52���4��%�9�!��OX���E]�.��mH��u^�Q9����0�}�&2U"�-�BN�Gk� -����y ��Zǋ�/ON���.��Z�@�ʺXW���ҹ��3��0>��:�O\��
~}g����ڿ�qP��2&k49q�x�m)p8�Ѓع�h�}Ub�Y�|Ȕ�wX�N�6�2��:ԃ�"W�S-�Kc
,(���5�t4Aj��E�4�s��iU�9�=�Y:%�t��s4�?/�*�k��~�_P'���RLڈԯ�RX�Ш:�s~ Wf�OG�+HF�/���Uh��B]��!U��`��\/Z���b�y�Ť���񥎝��{uf�-SH�<e}?������bȯ"�������z�iJ�p����(���y��#m���6s�z.���@ۃ/�#]�F'��`Aǜ�Tl��N�Tv�]u'�-�q����������_��\�>���ܺ� ��Eԝ._��,��o�<N^_j����D��w����\��`�U7�鐨a�8�#����g�A�v+���("z��w����۾/ć�y��E�t��/��s��Q� wq��uE�	��ώ�HV������¸��]a�� )���λ+����k�'����f��´m�~vλ������QB���Z���k�&�e�� ��kTHX�t���-������Dk���G�\��f׮��ź��a����IU��ǥ���T������ٌ�J����R��N�E����M�A���:����̠@�~gkB�'X�Oơuե]��xӊC�]u�5�`�l�
�(i�ݵ��Al��uĩGm#�|�R������4�g\'�:�rn~:� ����׺����6^
)q��oR>R@��]Ś�����#�?]��N��:s�Ѷ��{�|��}޿f8`��q�^�q��TP��e�M�x�;�I�P�9�Fؿ�������ɢ��D%D�uK���L	��`����˳*#�+Ӑ��3/�&���e�Qp��g�=t��
1��{��>ZV���������п�����I�ˑ��~��˛dTX8s�F�n߃ڸ�8l��4��Џ]��&qpRA�J��wD����
K�t���!�w�,ӎԱ��n.��zJ�=�i�
�%�c^�"ݧ�a-�v�k�O�`T�궷��9�j%�M^�eOq��[� �<�MT�-l��.֏�O��#"֜�3&�|��y������Z8f�譴�n����%�חD֧Z?z�x��A����_�]J��Xx��P�G㼟ԋ�D��N��cZ
k�d6��z꣖Av�E����)��IG:(�<��
�~��=?����i̠`��VC$�$DjB!룼o�Y��"��C����~�e�w��}�hv��(T����N�J�մu7Y��z��j�tZF>�`,'�,�9c��d�>�mڿR+y] �]��k���.O��5/n���[�v�����C0ռ.c��	_�dt+\
��x	�s]@� `U[_�ED��rVٝ'zX���� �������y��'������hv��������e>��:�i`'Dw���H�^�<�����l2�����e�/�������{�Y��	���<�+̋K�$+SX�C��b��:�,
��9���4�h<앝�SP����;�얈ڨ]�͓L�3�s�t�/z�Y F𠌶T�w��\�����U��C_y=민�f������ׇ��)���_�oֿY�}��K}�����=��0�I�:���
�	ඹI�l�{.̊��S��j{ڔ��Bo�z��w��ߛ����k���iwF��v	���V�<ș�y�{
�L|�^���.�_�&ޤ���Fw�����~9���ܴ{MK�0
���4%�]� H��:e��=SHT��GDy��QK{�ұ���1��/n�S�_p�n
�J��!�� ~]	��3���O��D6i�?Dw�d�=��;�^�:�;n<��b�I�3O�Ѱ����ڷN�?������n�i�ح�Hm�m��U�
�w)j����䱯�v�N8+3Ƶ-7[���U�E�K����v!���`e��S+��c5c�5�6Ųǃ�!9�Glt�GQ���E��g��k���S=_;�]���1��Sw�;w���Rv���A���Q��J����cMa��M��3�1���4��zZ.�/L�s*Ga�������i���<����:B֣s?��b�˄��\/��|B1���V�F����,�����:=�|@�KuM���	�����\����}y�D�	MIm���Y�7��M���`޷���|��wO��-D�8w�~j6��L�s��1�L�m�/���u��}�-Ʋm��[��4�@�R���N�~�X?��.�{^XM ύ����tl�_��g�'�,^�|PF�Hl1��/0WFx4ƥn�ל���^j��EB�{��xҢ^c4��v��f��=��j��)}s��Վ�6��@~h-����)˼�Z49�;к@��������MC�P[�>q�ʾ��t!S���|f[
�}_�� ����w��^���!���:��ܓglˑ��J����U�R��l����62β}Ln�&��?i��-L���/��y�lʦ�f�GԈ��%��*�J�\a�S-0�����|���vo�c?�a���*d��5#�O{s��1�i=���ӄ�^B१d%���1�+I��J���D�q�f8��RܙA��������=m�MA(��M����촜iB�yJ|Z4��"��e��֬L��bQ��I�,�I͵>JC�0q1Ġ'b0�r��1�m�Ww�Q��ګ�G��B��K�����g��5�`Aq�Vq�d����[1mtX�+�{���E���?��6'�u۸�.<^Ǳ�o������e������9ei�N��w�&X��e��-U�l��(��+��D�Vtn��a�>�8�}�Y����
�UIZ:|�m���.���	=j��Ғ�k
���19�u=�F�`���Y��E�z�ׄ8k�m/O7e��O������&���x:<��9�8^>��BwZ�8$�og��b��zپ1��O�A��i��m���[3l}�f��g����a�^Q��d1�t2S*Mإ$���k�X����g��jkꒅ=��S]?�����dRq���"$��tv�>Xh7��(G˼1��i_`�@"�K$_"-�N#�$P��ϧN��}�| ���т���=a�m���w1-��4� �鉟���v�m��!y��d�l�!�*߻e5��=�Ad#W�k82im.��s�r���&nE ו1l��zu�'��}�q���1��*I��.}�!��2o��\j���
�������В����<�Qot� ��%ѷ�ḯ�beʟjlk���:���s<+UK��S�����u�e�,���������B�av^�^i��7s������1��z֞�gt����u��lbpaUo������C�!�O��Y����!၎D�ZG�,ז&\�`a���(p�&���Q>�C�Vui6)�W�;E�T�Rb}���&�`�?��äv�}ϝ��F;'���=El-x|����#+��步�����!��D��밍'kߔ��6 ��%b�q͜�pՍ� ��J�"��B�v�|��3T�x���,�M<Tq���!Q�����4;6.V	���]�3������#�m�d�{�3�Y�7S\�b��'��s5\���L������"��wǶZ_�G���cL�sw����pk��>�nf��W��]륻�u'?��1�cD�.7��L�DS/�)�q�
<�C�/3$@���5G����r�T���fM�J�?�S��;)��t�k��I�.K�y']��;�����
&�7�@Y�ԗ�.9?4�wz\&���U�'xz����սX�,��<A�/mh5Z-���mR[I�&$�=����<��̖���,��C���_=*��|��CG:)v0o�^�/ǁV����^b�|�:,�ó�V�u���Y�����&��A���Ӷ���]>��H��u�m������N�h��$�[P�X��,�_�.�h�;E�z����}�_�M5�F��\�g��޿5���οf�<iq�F�V����l���z�ȸޘDK]��*%�#��Ȍ�F1_η����~�yx`
�<��R4��O��%H[��ڟ���B��&hu;�XPe��_��J��s���W֟%�[i	���n�C��xSs�D�W��h�dQ_���5�}�8�-�@3��R�]=�=��s&Yҟ��C?N���Z	��+�`i��r��!�!P�Qo_z�W��L�q�8�=7V�筓'	�m9�X�]Z�^|ڳ��Z(�)����ď�7���T�fX��*�J�)�� �aH���� �aV�.��h�r�m�mM1I髐e�c���ҡgLi\vh�&|b�q��]�Up���FA�7N��T��̵���}���T"竻�����cy�5n�L����4�������\���=�m�ӡ6�NF��b��W�c[���;��tވ��k�*/~X^-�ӳ��55������ҼC����ok\��V#�!:�+C���<5!���i3~�'Ĩ��@Qe}&N3f؊��^h��������xC�~�T��9�F��X�ϊ�{ӊ����9n_z��sN�N*�K����[��g��Cr]��W�U�'�}c��66����L�aE%dB�J��c�w��Hg�6�f�%�����(Qn�w:��d#5�g5Ĵ"H;=B�I1�|s�4
���0	w��nEyrm����`Hs�*�n�-RH�DLܺo�y�R�M��p�dv{�r�A�7�Z�ߥŴ��ݕ�L�8�|��`}���d�t��B���\�S����Z��V7����(t���4�?�6Ȃe���B���ծ��C������KA�C� �+�9�Ϟ�(k����Q��\=d��g��\��z3g��G��/K�"zC�ɸ�wq�z/����b�I�k�B�7���\����g�ab����Z��w��xM��է���K�?Y�t���mG�|.�ۥ?�^�
U�W�>֮,�{��`+��6�?�^� 5�j�k�����?~q���g��rI���'��$f��/��m��r��K�5o�\猫h�0;�	�|�����(�xxe��8:�=@��]\UБY���3�����5�^�����V�)�WF�_"'��Qȧ޻��=�cB+c�cm�XxY�n����:�Y�^af�t�| �j#���.z���[�W��O�z]h5尰�k�%仡՟ݪi�� {*C@D῞���ޔ��4��7i!�^A��s XM�S���?�4�ܲ�<��1�}�
5_u
@�e�dyG���8��+z���p[Ĕ���.(��T��L؃j�R��z-���G�~-E�i#V�̏תK@�P�/1��>�dwm��0Xއn�����՝,�/gꖶ��9�@��������)�}4����'Hv�u�Yv����Ϊ�u4�+����F=m/Yb��^�Lqv���}��Meb�{����-���
ʳ���E�x�6�������2��I���-��X�����|ML?����~�/����jJ�L�S�3We��3�@����H�)@�oX��/t����%�G�����Gd����xkw�:ݹ"^v�����$������^̀�X����r��$��ψ��\9��o��,!N�J��5��:c�;?:��8!Ѽ����\%�w�����A4�@(�h.��	��>Z<Ϣ��ŉ��,���_��P�R;':�Ӥ�@���cF<����j;;]}u�Io�-��ʳ�Qk�N�o7�v4�Pp�%>C#K �6c��r����s�-����t���'+� AC�q'�[N�E
�|�>���0%NOA�X�[���3�T�?Yj$��L����X�=�_����r��3ϵ�F6}мI=����>$��Ԟ���3<)3I�H�u㕑�������3���	d���B#5���������6�
&0�n\ �V��4B�/��?��DC=�����+̮C�Z��$��y��R��^���X'f&i���ZD��u��Y�N[��S�(w���]�k��z�3����p���ε���r�}���H�Ii4���IL���Q�y5V��7�]����M�� ��V��m��H��w׏�d���ឥf�Z0*�x��莅�`kg��DzᇲGWe�4:�2���;���ݑ�X[�%Y����̫�9UE4��[�ح�S6�T��ON@�u�b�x4Ѧ���Wf�@�,��#�W����)�[����r	SpB�l��!�he���_��qݽ2{km�mX�[�#�W���3�w��{�ӛ
��;��ҳ]0�Ա�j�oR�Z4�T>"sMn�N�l�Lv��3'9�e�_��=Dyѥɻ'�4�;�����E�9��[	c�S���#�0��R_E����~�K֞l�J���V�8m◚@�Eˆ�W��њ����@T��w6�D<�?�q��Ҧg�)C�+��F�|���5n�v?��P����F��D�HĠT�7o9,�#�rܺ"�-�E���]K%S�ڧp�&J�:*�ٶm|A�@���4����[x��\�Ygj��ݗ2��:���� YY�������.+�B^�������'(Hpu\ ����h�f\��
��p�'�/)�	�w���j����Rt�#�޶naY�t�m�re�����|6k���Z	���C�.X���!�q�$_	���9�R+�	�&"�8ƕ ��b��.o^�`�@`G�V��ha�,?Q+��x9}�k����pYn&�,E[c%.	K���d��)�<Z�^�"�E7���"�}�� �P,	lM���/�{+�V���}��:J#��z"��n�v	6��f%}5�=�k}�"6,��b<g"��U��8�nz�U3Z�y�	q_�w$�)��$I�%�=���+�g��zd/+�,���0"*��q�ʛ���w�씴4�+W� ��d��'���-XW�A�_�!�1�/�
����x�%q򓞳љ��[n;��\��zfd۟c~h�*R��N���Z����Ԋ ��NV�1�<K�	�;��ô�4x<�z �_>�B��cd(� c���8INk��5�6Z<�X.w$^��:�İ/���A�������N��%�B/矫Ul�%)+<n�4�
��&NL�ll2B�j5Z�^��k�\�S�����g=������ɉv����[��م�2�~�/λOK�ߗ�J3%!�e�Z3WT{�M`)�Mov9�(�*���H�d�n	ZP>���oc�����:*3s��|���VGo���|���	�p'QWY����ŋ%�_���#������,�-��]�R�l�~�E��L&�Zt'V�Io�U�"&b���6%�;� ���ɩ���7��B������{u�Z�O[�'���_F�vy�f�K���_Ӝ+_P��Xz�~�A�%�������2�$����'8
��o �?G�ͨ\�8���,����S�um4��D)��!��B��{�|������[�k��C´W�yю\���zt ���i�$CA�T������@�@���!V���䡺����V��:ӝ_\Ǿ*3`K���=+r9�g�ǧN��<��3Ԭ.{O-�dq��"^�����^����u�!9S�FIB�����:��vD�t������L�c,ˈ��_������`3�������|oP-~��0[����љ�����.�M^s�����4��nFq+�F�~�t�B�����{/8�K�"d�� *Y���D��C����i8Y�ϹMsᬨx���sr����B ��.�E�Zڅ���nk��y�NA��DC�]�3�e� $ëLT��[�yb���kPc��(~ѭ�Y�)!<G���B	d���2\UG�s�9�s��T���y7�.#�����������%�}�i��T�5�Ͼ���l���Ło.C����v�b��w�V"��9Hz��v�s۸B>����x�.n��?.9kj����=���3�W��S�&�W?��-|�$10s
%蕃m��gy/0,�o�|P��a�����v��_� ''���".�,��+!��Ͱ��ó�c�����3���)��wHL�jn IOvg��9�N�5��h^z�D�;���Tf�0�.}�ka��M&lP<�g���S�-���;<��eG���Ufo�ށ�0�D�\m����Q�Aur��r��ʝ�3��MuG<6�'z�S�R��\��[�5�Hf���#G�=;,�~ްPR�V;aۭ�S�I�I�}�B��S�e�2tj�2ؙM*7+�a:m*�@W���bۖT�w�Sb�Ɣ����q��{ʍ�*�	�/<
^ι�.����@t$�kڽG����14�B[	q3O�n��?�QZ��
�n��ܯV��R��;��/����C82^��.MEN�i�I�E�9.��'��gԡ|US_�8�
�w�X?��=��}��[��]đ�o!}�?[��~����W[?�:�r��].һ#�cu��-�f��*&$����>�>�d����f>���f�bE<f�I
��.`�'���� ���g����,t=�*ryL�9��R7�Q�j��8�Sߝf57&���z���O��f�"'���?�y&|ҊW��U�6�N,L�9���pJb�y�֐�%���?Ô�kv���t�|��>77�G�������],m�%�$�� �ȟ6�vӥ��)ޡ�OP�zVɁIo��E�)�W_i�H�2򣏩�@)��:�>s��y������1�L���ۏ��|��@x�����B���Mk:R�	�r3E/���\��Zw�������ۈ���n��H@Ѫ��֨ln:��fegΖ{s��C�~�¼sfE1���d�,����o��g����2`�H�\x��}��mc+B*�'�D{4d�s^'�8���7A5?[�+�|_���!�]G�}8{����§S?�m:�dSi�����v��f�h�wV�1\U������V�p�Ys�e+k�&�;!i�p}�,D\���n8p_Y��Ӆ.�pl��-0�t��J��[�́�=�`�����,�C]�";�%yuu�p��TgEV]F�G�հ��H'_mNE-��>�Y�G:1����~�[r�|3؛�A�`��钒`�2���7�����������ru�71	e�-�o�h�����r9;/�}N��q!���L�a��U��39T�� @�&���Sk��<�� 6�)��!�"d�j���6>��/mgsQ��]*�Iez�MlN��E�& �F��Q��{&E�nmJ�E�
�YvU�]��L�S���o̊��T=���<n>q ��
N����[�]�aN]��y�(��R���S�S��O-khwi:�v�T�g��g'���g +)�ƣ�q���&^��,wj�3�������ܲ�Ӻ^��*0[������+��n;�p�K���sL]<�ԖӢ	�;a$�*�n���Ȟ�vu���=��s̭|a�}�j"����އ�_���y@���B�5�Z���#&��%Ã\��T��6�%�ɯd%XuB�4�Ӥ���~�g���Y J���KH�{�j�n}\,U�X)`\g���d���Z���]^QAQ�-�տc����[Z���EJr���׮y���4�6�%|g�p�M{�ݔ�y'������i��,�Q�>b�N��Z�&���&�gѬSCJ�y�S(wP3d����E�%�وg���bԆ�������;��%Z��%�hNDSè�Z��H��'	�%5c�1���/��S�}Y ݐG� �c��v�݈I��1�6t[�h�%��Z�͹-EqC��vm�ra�H��Ojp��)S�V�!pR�6�N���cj��޷��'굽�I@Ϩ���.�J��}��Uf���k�F��J�}��)�G/K/�j*�OW��Sڻ�JH�q4H��T��i�'� ��� �㙼m��8���*�.5�{�:_�߈$8��`�ƪ��6X��.����@'Fv���A7x�������rg-u��\�j�c[DW��h�#cC�LV��ͩqhI;8��X�d!x ��A2�8*�����?E�'4�ǁ���J��j�!	Z���v�$�;���J;\:B��W�)�\�܆���gnSo̢���j�P,)��M��q�\o�9�blwo�۟E�N�ʏ�;��;\�b7�Q�?�z]&k��Y������)�ñ�uuTb��l��S����N�=�r�u:pL�I����ݮ<�._��R�)����m��o�sP���4��yt2qT�j:Obh:���I��dGƔ�[���t9,.�ͪ͝�Lo�T��q����M�F���5���=�a1�K�q�N&�+�f�:}ײ�����µ�HV��
9���"ȓ�d������s�XI�R?�������֓}��3G�3n���k��|����ReʻYw�b�r��fl�Z��Q�$D!�]��G�O1�,Y��xw��Հ��9�\�5��/�ػ ���Y�Iu��Ʃ)7UU�}k�S��Ѡ�n�>:B�Nd�����o�h�G�*3H��F�N�������|�*�y�w�����FjR�>�u9=Y�G�o<��qb�Ӥa�D`�dYx��V0�a�)��#���W�C��[j��jl@(�]�
��T��Z�N�X��� /y\dA#V�n��8}��
(����D�;��hE/��#nЭ��ɛ*�"�/s1�/_c�(v]�?��7���_�h��t6����`z~�fߎ{:�U�tag���s�E�m���Y[�7�E����_~+ٶ<��4�K�Q�u%h��VH3�@�S#v�a�����}/Ҷ(�K��Z�������mG`�K4꼔����+&�v&Qy�i��-LcIL�l�^Z�yZM'�����w�~p [���u":�O]A�x��QO���k��nօ7��&U���cM�f�Lu<c}c]�B鐘ji���5��L5yd!�1�N8]g�n}C����}NX%�Yi�|6+��h�_=��0�mgzkB�P\�b���h���M�
4�58nEU5ߤ*��p��}<�������2�(Ә��^kO:Н���g��vW�;�I�j����
n+�E�f[猗I@ׄ(�����6���*!W��3�e�n͋q�5f�t�.���%0��{Ά�!kQ�J��-�����	������E��J��)�!T+Z����� E�%E��V��S��������/%�&���լ-G����Cx��Ҋ@./Vv������*��T����9�;��1�i�6��G����I��pS��@5��sk@N)+-�,�ĭ��V��զ�:���x���K�C�g��2�5�6�K�+�M`�h}�P�K����ف�T�%֖�X�vo�]%#��:�mg
{3;��N�C�	����t�BQU��nW��G��k���g���������$-�O�j�?̌�!+6J�!�o�L�nzk��躰���/>�|ioz�f2���Z�y���s���rifQ��'���5�%p�W����e^�_����9I�֛���
#Dc����I@yM׎,�������������t� - ݹ��"�� ݽ�t�H7H�t�� ݰtw��._�<�>��ι�0w��n{�|�ˁoQ��w=�>^�ݰ_�SR�wU���f�)N��t_9���qʖ'�QU&��}ˠ}\���i5�Z�M�)^���tL3E/p����H�kJ���w���C��(f�8]���O�]	�}CM1m[ ��q[������&}�Fۃ>FBǻMQ�I X\Zw�Z���y�Mf��@+
ە�(���T���9�^�U��`!�M��Frcj�S1�§]�h�Z�C��Ϸ�\�4㿄Q�Մ)Q����.{�2,Ŀ���R�g�;7Uy/����y�.L�t�}�����?�N�n>xqX0����Ŵ���L�X����:#j��i�&���5���'|�{f]b���6��>��0!�]\�\�>
A���)H�ћ;����W"���փ�M�e��ބ}z�K�����09j�l9=��3U���"#%���t�p\�DG���C�Ƿf�,����z��R�����l�xRY�ds%�`�w��32g.�y��FԚ~�B&���;�Y�yF�.cӕ�KGOT�K^�ڳ���T���Q���N���}�v>_n�8-=�2~YY�*���+M�絛s�.
#q���se��2v� II�f��b�
���Tp�����`hQ��՝��e�cI�I��/a��D*��<����PO�p���d簵��7�TB�F��CR8�k�ŸC{W�� ��(m���Xxg�2c����3���"=�@�֔eD)OI�x�ʦ�֖�x�j��I�vc�!Ԗ��5ugT	�����
&��O�ug@��=Y�eC��m�zH��{��iB���K+,§?���9A�;�=���z��~ꀂ��iTԍ��y��T�,��Fa����0�^�9m��r��Z���<��\3�;�xo����K���8|�╺7��"W޹�d��ڥ!=X��+b#�W��+Ⓝ]|h��rX��e�"�=��#�Q8�i]5t9����o����J�䷱l.&1E�WG�`�r���S���}cȭ`��m�u�W�B7@�E�6%j�~�a�fpm� U�9�Di.-���ˤ.�q(O7�#��fjzM����#A��R7�'���?��D6Q�Z�5X�t6�@-�I������ɕ	�)Q�co7��e��r��
)�	�JI��O!5iu~��S��w��ѱ�*xQj7�)�?��U�o�Yڳ҃d�\ƒ2�w��&5U�L�IY_T�B�uxx��2<�dv��}��&'��q����0����D�p9v����^>35�s�{�������Ǫ,�$��b�WZ!���Z�)d-��V�;���JW�O�+�+��Rb$6*>T���no�������o���5cHCZ�3 �>�<JF'�oy����z$V�WJ��D��@���T���L��
�[��2���p�P>W��:~�'�T��TM����d���jVs���vJ��T1���\ݛY��CǛl����;�j6� +7`n]H�]���a^6ϯn���v�PZQ��cœ�~x[t����E �f4��z�dUۂ���EU����Nې��F/.%���S�����U���K��U��0��ġ=t�f�֚I��[���l7�^'m�'-�5�"�$zZh���c��Fi��!M&�1L΋Y�ȯ+�#��Ml##�FRko��&ص�ԃE�)��N��ͭ{IS(q/���>����!�W]͆7�~��O*|;:6:�ܥ����]pHTvH��/�zh������J�	˯=�N���D��N|V�R}�f�J�Z:����fW��[��*�F�S���kw�yx�/�&\7.ə�p>ю!;o�W�U`��K�7�<��瘯u��.�d���P���3f�Gb��r����(�vw$j�s�S��WݖtrY\dK�c9�=]��" ��`�n�7���:*�R�7x�1ӏwV�=_�&�M"
�����+ҢT�h<k߂�q��Gb!�#��P���K]U���AÄ���:9Mǈȭo�T����Ԥ��Q�߶-�Kn���Ro]��\�
�Í̌�b��&ˮ�����w��z�ZY���X>:Q�Ⰰfw�XϝnUÉW��NA:��Ǚ:X��JXH�7����(�bWU�ά��OF��T�葵� |"��vA,O�K4=��F�$w��SIH,��7�H[bo|Z�~^h+�H�UM��P)s3(�j\�B�U��o!g��HQ�h>0%+d�X�_���bR��0ӽfl䴏��dV�pρ����p�9�-q�$)V.sr}A��r�)A�׶�qJ􌠡o�>
!�{�'uA"�=(b��]-#��)�Q�^���c0�����D\h���hu����eƘo{ת��ڷzC���V�RH�&�R�5����IT��u>��r�� ��_t%����iզ�ˌ�UX'q�4��yQ���
V)��?�Ü��-W�|�Z�	��X>١�D�0����p����2�TmX��Xq�<�BO�nW[4��m{8�}7m��^�F-82^����3���FҢ�]�γ8rl��kMI�(�{�,�]�rNvY����[��$W��=�>>A�<Êvj�t^�N-~�Č���K�tM��1c�oA�4w#|�w�}�S�`��=�:@2�;�����7\ҍ���D�{s݃�T�1e%�ջ*��+k6�m&��G�*�ɞ�|"nǢ�4y	���a�>���~}��C�F$����m�p�d'�|��fP�V��+E�'r�����r�߬�B�JRP�YgS`Sn�%.�8m��g�[prP�0bJ�����״��������TY���ay[u�X�^۷�W����)R��l����~���~����cx]�E�bn�Osj	E��$��4]�ct��;����	��#����Ȼ��42�W��ڥ`����� ��,�S73m����-2 �L�z�>��4؛�J��t7�uy�t~�C&��+���T������|7�,��n�U#����.x��Q�d�?;�5��n��$F��'�0Ԛē�:��_�JAUڒz��b�ױ�������`�S��RH�3���١�L����o5�UC���]�����ާ'�ё`J�s>w���*~�� ��V`�
��A��M�잸~ѽ=]�v���P�ű~ܳ�j5�F�����c�H�Q���=����כs�Y���}4�l��Z�1R�{���:ͨ=N,~���\�`V �\�����<N�����>3�IpeFX�{��d�֍ϧ�!]��m_ޙ��?��r�]r5Վ�Y���-��$������΅�����`��ڞ�u�T=�y7y���x<!vjbU�\��~�B���{v��=��-� 7v͸noS����QD?mo��J�E�&t\����ʏ�N�����a���;��݀ݕ�k�E�ɉ�˰?'0�	��&�sD��qZ�Q�0g��ڭ�T�j�OD31�p�2l]�:�#7��d_۬lB7�+��rs�4D�m��R["�Z]�A�5R�w�N�jH�飱R���7�[+O�Mz�oC��	�
�1|s�	���b����eS=���;�s���L�&���H(��k��ڬ��;�+_)K��}����W'0ae���9kp�_�(��$=!���0Y$t�դBT�����x�]u�g)�9��t��2p#koAC-�� ���*�׃��/4�,P���p �ݶ�	M�m;���6I	��>/(,/�c�Pͷ��A���PJ�Phc�N��w�-kݞ�A+,�SL�7 �-�V�u���@�Z�9n�fH�W�.�PE*�����޵i5�_�3���i���J�2S3H�b>y"���~����As������[������&d@�
|W�C�~��H���>�n��ڣ�Zbw҉ �~K�FB�$|>�'�@�����M���߹Ѩ-�qwE����敱�����ꨶGa�|�a���u{��Ǌ(��S�%#p��F_"-�>�|Q�`ց=�=�&È���s�<�#�j"u)�)�
��s�ķꐍ:�C��dg$O�d��|��H���Ŭx�[Q�S�/���D��.�NG�U�3®g����}��
��l5S��9�'��njZӧ���U�x9�q3�ð�K'������._s}�Я�o��[���q%�*�8]5�bD�
c����IFk��h
�xY_퀘�,E��ɷ�D��|�l�-=<+`p�+�̸[��FkXc|q�zwsR6|}����A�k\�����=36��+�!6��dn���F�{�|���02�xL�4��៷�;��A�䨤y����8��}ٷv�<���M����譅�V�̩�Ŭ������~�p\�p���'S��g���pd(�5A��V��4יJ���lipr�=R�z�l����U�O@�WOdk�k~s���M(�n��fx@�\[r;
�žU�~t���������_}	�<��J�r����W(��nai��̎V���1�"./�r��gk�\�l���lJ߃;�[�ikE3���9�"������=�3��2��s�@��-.�x�2�K�d��w�iA5�}R�y������a?�\���s��	߲�_���@o@&�W
c��G�Y%��A�`�����M�Z+��'� �z�9K���g��C�,R�����{=����Dd���0�<~�;:OF��?/�#l�X�
��O=U�L-]��!��E�|c��gXݢY���0��G�~���1e���C��ޜO���	9 ���@��`�7Q���-�%��f;��3�+�͵ͺ黄�.n�;��Z�k���s�D���-n�/�яz�Ff�Q�$F�����L�T�/G�b����>���ĵ�k@��z9_���㍥�f��u�����6]�\Se�c��fz��4ʂ���.�_��3ͳl�O��U���W�1�	Y��Ь�6�6ˍH�����V���&~�G�N��8&��r>l@]׺�p����[���e�}7&�d�@�&='��4��$��l�C!x���~�϶ ��Rs���d�b�2;�.bl�H S;QIIFS\�ko�(�+Z�l���4�t�q�Ϗr�#A2�1�'���a@ZS���=�3����:>m �?�'��I"��H�����v���?�J۲�Ү4TW�m�78u�N@XS��v�[S�~kY9\��lp��F�����U#�K�۴A�6��1P,
U���h�^��Y�r��/� `��"(@���xW$Lh_��K~cDi��F�v΍��>��pD�����L��)+ȝ�*���]BY�1IS���~j�'u/�XA\6-�Pi\��r��^��9#,q�-/4r�rp1jKe�0^J�����qT2�
� �Hu'��*��C/�RÕ���� o�3���s`?`���-;�(�Ȭ6x����(�[��"�̘~���q�u.+�rf�D��"���mqN)K�nyS�`��G}�7��e���	��m 1���G*�Mg��aM���f���k�3ML�ey���QP�z�#1���ǂud���@�ɨٞ�=���v�j�RҌ�x�WT���R�t�UX��8PL��`h�dj+G8�_��yJ�l���r2u$=y�����3�>�*M�ʬdV�M.nX{���j�]H�6�e��i�t�>�����7��:"�(�\�۫��ZI�!�@�8�!!J��TM̯��3Z��
gؤj����O2Z}�Z[v�KRBw�G2���D�=�-��U�+��@�7�sv�Ǭ�\˖[sQw�����4竞0��;���=����[�/��KL{p�=�#����� rb��0�8��`�A���I�Y��R���� v_���x.�K)6��Melќ~#* V$�ȟ�m���-����l�gU�/K$[�D�0u/!�
V���"k��tБΰ]�%�gʙ���v�g���]���;\4��^�.~:�uh1��$^���޷���7��k��$a1\��������%;&1�����:Q�
�<1�X��ۭ�K_S�L!��˿��񄊜k{k�̟��<�wh�K�ug*��pk����N�LD����P�I���� �W���l>�\�2���^$p�5����7B�.�`U��:LD |r��cft�saK5n���-h��k�y�����c�-�,nv�$ef�<�2��Rz��T��}?3�??��|N�2�qUI�������CJv��s��ᆓi&T"��J ��,we�}���L�)����tA����IR������������v� ���^7&;$��V�̡��& m��S_�����c3[{^�g���Q�h�2��Zg"7n�_̻\|�k�½/dO�t/�/2~o��W�v���ƌ��Qwo3F,��g�k	l� ˠ���QD\�������%�������4�<�l9F��yP�M��,�"���fa������vq�f�͒1M۶&A����.?f�֝`�=E-a�����E�P���X���	\��{7�� ����X%�^~��[9��	��C��K,J�0ܾ�&��*M��^���Hב`��T�dZ	ѓ��2�S����w��a4[Wb��k��k�u:w����g<���\��	v��k�^Q���T	/�ϙ�ݖzU�+�p���aW.�`�QP��e=���h�\dD��/=�9�������R�P��ӊ���A�8x� ��}d\�ՂHo��W��8�f����&�r�F?���λ�;�EF��f�ظ�_��&m�2���<�#^�q֎]�l�q����}K�مA�*%bw��֓��w0�-q�T+u��{��طp�J�ϯ+���}	��
t=v7Y�9�@�&�@Jh�S���:��*b�{�nv��PS���Y�І�ڕ�sٗ:Ɇ�Aa!�Z�K�ŦlW`��~��\ޚ�'\k$�ͩ���9��{�����~ċbU��ŷ&h�C�EO�R�y�Rs��d�����S���鉮C>�n�#뺞��_NG�P�Ҩ�U�l�+�r���H�_�؃���=`}�@�>;�TZ�o��r�e��Y_9�����*��g�t��p��:��(�ؼ��CI�O�-ߏW��lN9���|�Ao΁��ē�|x4W��%o������m����-�.�zS�ˬo�m����y�"@����z<�3�羚�`}����J�\���)�ff��N��82��i�ms���B�s�a�f�t�F�b�Ma{�|Ç���cWD���F��}*���1�u��7B���MV"� ���5��u>�<���)W2o�sn�"�P�����x2���YF��>�;u�e���9l�pHH���z��By�w�H�uA�wDx\���#��ӳ_���ZWfp�~��%��%[�V�V��&X(SL���{��K���.����#����ZJ��{����}���'��Nw5	H��duM_� �}_+��׬u*8+�A�A^sn��)R%֘�_��}��^���0������WB� ��`r��<���b��W��>(u�k̽h3:��Ƿ$9�:h���N7ᤦ�\n��ߋ�c�]�'hO����SB�v�x��[�L�j�]��%5aq�3p2������By���U��u���wj��/�F�I!� �qf'�݃ܤ_��II"��Թ�`k�v���a�(�y涆��@{i��T�Օ��?u7�vϙ3"�<����c�d���>"��#Zuut �\��Y�Q��4�Y��?�'�x]vk"�m6k�S*;�[���Ļ'~v�%�<�J�f�A۲I��(x�3��56��:�9�vt��{z��.+o75
���y�͙�yW�8��z��V><z���jY.���O�;�87:����jxͽ�R��R�P���zc���r�z���'��n�&�`Ҟ� �s�=���=:[ѽI|���jYw��p�	�ep�5�K8�����Q�����+2�f!�������D�'ܶ�PN[��D��0+�O	X����Q�R��o�d��T��w*J��������v�AY=C�j�K��`5~��Cm��&2"�����g���u���
ߊ�Źw�X>��_�p��K+{i|���{���w&���dc�Oo�z��ْ]�wvZW/5c�=d���Z^C����}{}���w��(OC��֍�4�~�hՎP2���<@9:�����F�?����w�I\~���)��/p�+��H׫���pCZy?8��e�&<e��Shh��ܺ�I<&M�|m�=���E/�O2�
4m��c1�q����j�����ؙש���գ��,%�bځB�bt�ޭ�m���}���V�k���j��m�-�'0gٻ�MZ1�,�ڒ���Ҧ�*|
�'����1��A�/��c���j�c�-���iz�\z��h�K�ª��K�"3o/Q��z��hk���+_���4��-��Q�̪���j@0<ُu�K����Ƿy�JJ��KֿV�5�+PH��s5��y�=����gΘwz�kSjC1N�RӦ'7��(z�/c��T{�*DN�rr�� �z׌���K@�M�e�bbqf�ã���SWzi��Qf���4�B��Gy����hq��M�@j�Ms�qe��|���?ߪ����o?̹�:�kV�Yt��۫��N	�٧�'�i�Tsw�Ҩ٧�\���p�5�h�H)��:�Įt�*=NN��)p�"[���!_+�AK�W3�f��QG����s��֟����@����~��%l�O��'%{Ӿ��!��s�·`,�r�Y���}��\|A@�|��c�M�y�ڮgY�&��M��_�߰�}h�0&��j|D��Vc�*&&(^5i�-]nע�ҭ�$6��(�^)�����Ą���L�Э��C�[����;�Η�dϙiS$�%[9�K�J�~F�L	$"2�tp��H����EZy?$�V݂oa�^9
�� Ix�Z&���T0��� �y�/�x?��p�)�]��.�t�=x��\i��a�YV" O؝�.gf�@��}L�m�9 .�Y�������\����m�Su�J�w��Y�mdm߾/m�/���(l�V`�J�q�^��7C������t��[7�(�f� X>у��^L�E�ɏ����'Ad�>�"���c6��S(wY���&���3Ö���%��M�%������7$|�1$�:1ּ�E
jO#0�����d��rt�P�OS�6od���G��l���d�*2���ZN�-7o�B�N?M���ca�ߵ�2X߯)ǎ�he�����"%}��N�ď�_�d�[�V����z�i{٩h�h�L4eD����m�A�[	���WpQ��XGo`�>89�[�}B�O�H����<��<-���S���b;�}m�=do�Q�����Ef��|�ݔ��Fw˭���&$!A`U]4���$�B�XSOY�"U�o[�%:$�Sa�?�e4�=��BY�Lmh:��
];�?��<8�9���Yj���<G�nG�0���j)ω�A!�beA��x�#���[�ߔP����Y�,e��k"k���f���V�j-|�a&�:ҽ������J�D�����"qP���O�F��"��'���&N�u�0@,��.x�����ƨ�N[9�}���w��p|��|��j;�2�S��?̛|���Y�S�p�]�E%v������.�O�O���ǳ'b��� K��v<1�$D�|�F)�&Q��,\�G����|�{���l,�'{�������d,(��F���3ɓ��6�V�E
*P��R`�w_�]vE:�A�]1i	s��/ar��#{c�����z���fK���D���y@�	�!7T|�H�6�:�"b���t^���0>�,gY_�LnڲI%|Č��������6Y�LR:��Np*Ţ;��I>�l^�A�/���1���N�x��ݣ�K1;����m��{
�H��TĨ���}�,q�W�I �sQ?v��"���v�X�xG�*5E�0�~2?<�ʶ��|��W���CD�/ßu�~�Vs���9~��������7�0���+)�������Dx�W���p���Iy^���:�R����`�r��_R$�#N���-z��ц�H�\k�� Rh)
:	��;^��z2HYHDD�������ES��8���*�笉�k����#tle&Q
�_uA����ٶ:6#�񾇬�w���[AJ��/[@��P9�M󢠱�H�rd)�V� C)J�<�Q"_/�7�̋2^�_%&���\�����ÿ�lv�Jvl�ӑ�L^�;dΪ�[���j�/8���?ޚ��sw �����7h`yG��K}�
�O�����w��RJ��f���̯��hj..�jf�az�TVz>�y��Dgp��F�Z=�զ�0���`�x�?��Z��?�nwS��S�pD��.m,�lzD�\{����פ���&�[Ë8(1ȶKhg�h�����;��ٱ���;P�>w�
��o|�9@����Do����

�rx�E�_8����[�#��8�p*��<�vxb�?w+�(���Z�d�A�X����5���!,aa����HR���2(P�R(f��&�����OO��ݕ�FQ�)�~����\�����'$�q��\Y�
Ȗ�0~\5ͯ�$���u=�ζ��N=l�O�T߿��-��=i����r��%Կ�b�W�҉L�r������+����j�]����E�c�>1D�s�#����E\�yX�&5&����&�m��8,@��K����L���?���+�ڀ��V�GF,[��QADB���z�I̟�}ù^�n�7l)�����ǀ�z����b-90�j�J�jE~�;J�Ff[
�7=�[�H����ރ��9z����Gu�ǭ�~g�p8m� ���]�ё�V�#Q��8�@�Խ�7���.4��O)���?������"��X@�d�%=��D������`��ZwW�V��z(}$��0?\~O�?�|�4l_�3�>��ٜ~����C�Z�؞�d1r����r�Oa�؛��w~�nu` D8����2d��6��L,��~��Kء��Ygfj��'C��_��S�*>�߶������zl���ް\	b�F����.�!w��Ĉ�_��b�}m��2>�~�[dU�j��N/�?��Ό���F�ׇ�.�W�j_��,�.#&�1��]A-�^�u1���MMt�(��B��P�s����@����d��lu�n:6*m������P4��g��7m�X��e;8�b8�?32A�w,r���(ž�����x�|���3D��*6����d��%�*`p$5J�\�vP�;�CZQ��= �=��*+��Rw��� �;���~Lۉ���7�.kZ�YA7�9�A���ͮC�����@9���jU����Υ����f���C}��Ugo0a����ۦE�J{U���mj�V�m�t^U��pp$�ϱd�}���s<��;k�
�A@�\����rr0���
���Ev���b:*��5x�v|��`H�=j���'�!�T��?�R&/2�;��ӻ��\:͠=,!�e�&[!��]��@J�7u��Ɖ	,���]�c��rL4���_��h���x0�EƂ`�~}͈(d��8!4]�T�|���h�'���(+I����/���LU�_"���)�
���=O@Bby�	Y�a�� � MզA�qa1����{~�X�.�9¯�S�6ڤ1���(t����`��D�{����ƧW����)�I�K{��2��Υ�%�'��D�A���fq�cgD���g%����G�:5>�`�T���EdYS�����Wj�� �R�˫�jS�� �s�#��^V9�(thi�(����(FI��~���t[(�f�D-�{�V��Qe6)��>��ih+���\�ww��Z^����d���xߑ��|j����u�����bi�pSf��[���@���el~-�����2�̄\�<��Ie)\ �S8M�WC�fC���;�ĸj��?�����ѱ�����7��	�NE��@��"��y��v�B=�$	���� ��5��{�Kv��c��܄����v4�ߵ�ټ%��P�{���.HR�l cc�C0�]�(6Km������<��Whr�{��%�ۨN[�AEQ�]��e���_�}1i, �������,32=�+l�EOc<����_ڈ6%�H)D�X���A���L��?��w�S`��*�������y����v��0���],�Y�4��y� ��$R��(�������p?-ţ��5xa!2�u�/�*�m��Ve�WO�q��=�6�_�W�^��`�� ��C��_j�� �����7B���������%���2�4��2Ѻ��*e 'J����&�.}%rъ�n�]��>p�B����r��>�Κ�� "��(�|}D����w��������l���?���l�A$�L4`�6� �(���SW�y��^�����R]��ڛN����X�T���/c7����Uܭ���>}~=q��ֶܿ��F�����P��N�W��ҩ#q�*Luq�����[���Z�y�`ǥ����Xo +�ʍ��W���O��qfQ�=\�ˋ\Ә��k�.M��kӇ�=1�@�)�8��E}�o�T�����b�����tN֍����8>d�XrB	�HH�_ 
L\}ٹ�Ae��*�%���	�z�k�_�.D�J����þ�����	�4QA��q�D
�ۥ��F�vϖ��u+
��q?(ö��h�3����ז4��z�F���9����x�|�5O��G�Gz�и�~�����p�*��`�@e��љ4tJA$\ԏ��y�[s�F��G"���~�:j�,�.8G�M�x@�=��y�z��
Ĉǥ��Mf��}2�8.�T�Ӫ�����������t�1֮��G�~�Oond�_�������hd���Eov��E5 �uu�~m��O��;���3&;��Y	����\�{�c�I	]L����%B Ic;��D5�{@�.Y�;�^.��&�b���{���{�Io�px�pK���v�_�R��TUT�'Ar�����q	\�u���J���@OMs���nّn�lX�L���V7��e��`��D�M�G��:(5�t[U흻�gi����W)��%/���m�C��eW=�b/���G�#�B���֥�~��o�ם�~�MR��)��e�y��"����A%�A�<u�)�@��9�t��&{*Zױ{�oC�J���L��"!t��%����9���<��^��L&E%�X����~-��+����4`�WMo�|��śf+�ot�l	8{��F�aVR:�s�#o����?�$��X�7Αh:��@T�gTW���%�0���Q�T�x5��*SMaD�^�'�����[�;�`6�=��^6�mb
�;�;���a"0���/�����5Is9avr��~��6���}6m{-�ݏ����y��@��!�q�s�%a)��kט_/�3�:g_�R܄�[(�t��	�����|��|W�"���}nC�1
�	t��9Lm�q,Kj�Xi���������n��kyO���,�;[���O�.�.и��J?�`�)#{kr���2�� <�o�F�N*�}�c�9�ح�(>#O(�lk�#�n�����*]�ȃ4f[��H��c�"���gR�l���rt�O�R5<L��%Z�Hd��*�����+���o,�e��*[�Ta>�����~�m�ƍ���J9����uC)����Kk
��@�j�e}��?�r��+�-K'���C���h�k^���'�<�u~�(�IZ���n���@} �����C�~#�S���ac��	����&���z7�c��w���WNuՎ9��08��7��{o�U�;�I�0���_��G�<���<�����n�\���B	ԭQ��k���4��,/��w}H���Xۋ��X�� ڝ� �֙U�qq �}�=��`hqê����Վ���7| ���5�v�QB�l�E��ڋ<Uԥ�`D�&	q�˳Hg7h���K����;0�9r����~��Z�:��][�k��Mg��4�o
�)}�q�N[c��޹�D�Qrq�Uӑ�/e`�p��򸈹kޟ�����}$�A�
l?g�h׽S��o��~�t�n�3_H��p��Pq�sl�G��wY�`Cr���+I�p׹��9��-!0,:�j���ci���iq��~u}<�J�n"�:Z�Pt@m�҈i54�NӢ}����+�Ѯb�՟I��5��%6g/�7v�+Bx%){3V$�D.a�~�O�7I��D����Fq(�
�� 
eЍzPyuǣ���29�f��P�J	�� �ܗi�y�۟/r��5�i=Ј��h����� ��P� �X� O���g���c�hLĆd�GB�*�c*�5-U�0�]S�ATdB�U�,����h�v��D��u�/䬺���A�6gw	R�u�3]� x�9��Ad��n?6_�6k��v�wەI���w�#�j�A�~���~��%��՛�!�q����;����'!�_�ܲ�o`���}.�G���tt&���.'���68�6jo!<�2�5>F)
��z[I�]��x�	-��x�jK���"|0�D,?0M~�/��ϙ�5��Z�ۊ!�?o&F�æX�0(��Эo	���ە����X����9(�ȿ�b�G��;(�F��8Uq�#�@֚�E������Rl%��BLlXJ�4�)ġ��T	�]��dL���3FX����MڧKP �Σ�@'��2����@�sKd����܈��egMs�fMJ.^p����ݓ�JE�`hk��we�2�"��*�3�N��/M��R�&����m$x�����<���ʊ��et�������&�#�P�Q?���Ɵ
�y���I\��0n$�첞��s�����ic`ˢ��>s��u�,2.�����b���/(�Σ6��Y�߉�Ui<�k��S�\�Z6�k}n�[,+�x=WL@5��v�(yl���ˏ����[�Tv�Ͱ%٢oѮ��&֮����i���Q1�5�QR[�h��k��ξ�A�>��v���cI��M^U�oGD���4�m�#�*��\�FHQ?�DoJȑ/]�}��������:�f��AC[�q��X߳=+���[��8�����:A�#��iGvMR:D���O]����_*�𑇀�DX�v>~�����VU/ik��v��~b[P����wgf�D����ts&��c�c�+1���r[˰�N��?/�	��k�3)�2�?�M��d�������/�-?�>����Z����#3s���h�#`?o�쑓[?�oc��e�$m{�6�0!��oN�Кs����C��%���0� �ᦜj�wb�!r)&���Č���2ug�J8�wO�#a�X�~YK�1�M�����"��e��çem�MUt����9}g0�&[2��Ԩ��|ܚ��wN�A�����Q=ʳ�NR�.���آC?�I�Dwt�iV�7��cL.���b��z���7'��%V�m-N�oT�,qv�&���[�zL9��K�qsuG�}��\�Gl��ꬓ�m��So�k����M�+6�H"��.���,��$���@�;#d ��5�S�-���:���\����DV|��$JU�3����3X��Ԉ��vw?=��"2{˸�d8�PuM\u��$��ȥ�0ob1��Q�x��Li���ԁ�����i�&B/�}Mmm�ZSz���0⭍���*�r�Ɂ�"���M �����? �Xv6D�o�z�Yo�����TL�#����Y�l0�Z�#��%7�ƫ����͢�8�����7< P��<�?��z�2�,
\H�w�����V:�%�c���>h��T�Z?�tF1)�@�s<���h�ƻN�$�us��ncT��zHo}Pp���D�	�z��������h_�.7��u�/;<�_��Q �Q�^���d]�a���Z���$l�FM(�5���K��-�S������������;����^�0_�6W�����������S������K�f�IԆ�L���ڬ��^Ï�:i΁)NB�tM͘�X�[yQ�0���)���WV�d�8��`L����ȥ�t�c��x��赵~X"3�&�fn��*m��n]L��Ɋ�c�N%�)H�lg�xw��ϖjTe���?�ę�>�wŭ�*B�RyO�X�N�{�3���Q���� �(�+UI����z����vUk�����ؙJf��XO�ƕ��{=�0R@�!��L5�@�M��9��&9{w~����?}�#����8;t�@F�E&�|ּ���K�9<'U�Ci^���/v�OR�vY��@+�N���6<���N�D(�'~#h�k����E�G[�����7pb�����0�����������k��XpZ��L�'�q��
���U|���В�R���b�Y��c�@/�r��'��v��kp$E����dj�5�� ?�2R��dKT�aAG������Sݒ��. >o��Зe�?��9���Y�mۚضm۶m{bg��ض&v2�mk��o?�y����k�u]��꽺��Vi1&��%!�7QT�Ao+\O���/U�z]q�oW��`��ED�S�TWkNa�d�X
YQ��!4�K�m��'A�f���}�!��ĎE���Ʊ��q�2F͵��8�S�����D��@3�y­�h��el�b���萹����0Li����N��P˰��r�$��r��o�/	OKg��1�� �Ѡ��o�j:VX�µ�K��	ξW!�'�7*o68*n6��贮j:Ɏ�N\:��%t�{mC���`7cXa���n�K	=�7�H*�#�"�P�t�֘{��xR�dg_e�i�\̚v��#x/ZO&�#�=I���xZ���V�ߕɶ��|����`2B�ED24}e]��j&)�5�E�I:�	�xj�� �\�����cՓx��j��� �;wҚb%	��yn7i�o7��S�C\�Đ"6'0�6�|��x���M#M�C��c~g�ݐ�W�vS%(b<����]Ep��Ph	wg��0���AZX�3�U{��i;�]���1?�~�םA��Z��A�(�"~�T�n���gʤ0��럎_�I���������X�c��.n���>���\���/�d��x��s5���
��ԛ o��?�7&[$��e��Ms#6�R�����/h	s6$S?��U��Ri*���,Ïp�%-�a=��@O���v�ݾ�@x��]�rbͻx�&�9��_�!��&u�-�40@Y� #��j�e��bP��>��&�b��bAF%��bT>=2���:����	n�$wH��,�ԏ��
d���G�U�މ����݇�!�%R��ˆw���槷
:
E�|�}��H�F��\ x~pdO!lCwn{b��g6#������J�(�-N���.�-A_��}f�'W�K�7uB�s��e�����Z s���5I�`7Y1ں����0�Ըct��s�|N��}�2��$S6�d���߿����k'����vR廞\�I��r�}��7�O� t���������A���鋚�`
�z����4J��q]�n�)7dTE��9�s¯�A�E��\������%h�6 �?�?~^���&��ėIWGy�(�q�����c�L������;�o�R���ڈc���J]�/!��$�F��z�z�~���l��i:��$m��3:N3��-�!?�����X�6V�u L_�X�e;������1�_�M�n��#�P[O#���R�9��]iЂ'���zx)���ћ`�+�����#���'���DM,��x7u�ې:7���~Ժ� ����Y���Y�]�ޔ?����YrX��$M���F�P̭���!��-	|���E��� �I���kcq?!�1v{WA��pI���+$w�Ң�Ug1�&���g��?��Zu��/	����<��x�w��l�W��Q/X*�>�R����??FV<�B�1�jA `� �z�k���GV�TBKR��Ō����{T�'�ڏH%���,G�	f{j��%F�����t������_�'�4���n�i�< �Z������Hy4��c� )&�,`ʡ�����q�l�E/�PEa@A�K�z�Lv����<�I�%!T��~��^G�gG��;�J�A䐣�\-Q�=X]�D��L N`��Y^�J';y�+�������J��s�kh;ke�Q��Ş�͆������Eߚ����s̜�莲^�:��vWvWBXu��_��z����<���]��.�*�\ږy$y���(h�H�qb�(�c��ƹ�c<�� ����>�'#|W2�A0KZl�;2�8l7(E@S�	>T��uSm���& փy5R{
�%d���<N�ɑ�!z}�]%��q
kf��C|�Ą@�! �4>��E�e��DBCUw�o���1lK��oZ�{��
V�ޚ���4�ط�0S�k'9K�B���O����)��������o�w�$��L=`�E|Bkā�F�0�AL���rh	��xI�GT��r���p��W���p%?�k��PU�B����M���ӌX
��6#(��(���l��+�L�K�v�0��^r#@V��J2S&�(O�9'��(���4~��{yχ�4?�
�z|7̓���>�4�:Iֱ	Ĝ�ӷ��v�H��]v6J<)}C���oH�!�~�0���o��!l�ԑ�|;i�mI�c�F�I9S�K�����6��йq�љ�)��љ�\l G+��-:��7_xk�� \�q���)�Zbұ�N�Ҡ��9J{kpy@ 3�0���~�S�\?�# t3�jb���k+��脛�=�.�/9�,�5�a8�,�@�UR4��8o�֔��+��[�z�HhR�5S��9,�#{ ��DڸFQ4�Lk�-����<؅��Ǎ�D_}V�>��f1�!��P�+A�}���9j��{^o��V������#�c��5ˬ��dG&�A@[���Ȥ��P�wn�B�$����w��"�6e�Iy�"�.���~a����"ZiM��N:t��8�F��l`C.l��t��`�n���ֻdfV��y����#�
=&b���&�L��>t�	qi�'���Q�=���G���ke{�V��e�M�%�����b� z�>�?�D��;bfOR>��G�^��g����F�؟��#
0��A `Q0Aڍ�]�����I������fe&�Kr�U*x5}�75���x��T����6(�D�PW<�2�Bx��7��8tntu�l������BA�D�K����s��*�,�wg�����®��L"��gLs@��*iWctIՍ��`[��ѕ�߱6�fm@p����3�X\R�����,�'ux�X$Ԩ�̟k>b�֭�������f-��&�W�EZմ	|9�����juM'3��}q�Y��r�q�MG��U��k�ub��C����1�Q"06M�*�<��۶�U�wL̴C��qͿ��\,��\b�"]�}���k������h���$BA�
cg�	��e;V�Ad谻iF�y�{��(��m| ���*�"Ñ�|��)�!Q�������)���f24>=L�� 8���k���V�d}<��]}V��eD�S��/����`h8�b�D��Ƈ�����Cʒ�Ɉ��T�s!c�qvQ�y}�sJR��L]y(�/�l2:pǽ�JNf''�m�^�E ��hD�y)��/���]�B@�	d|�41c�Gv~B(�Ƞ-9�ر�».��VЌ�� �o��#R0k����Wǣڝo�ˎ�H��T#8�l�ӳ��ZB!x�����8��8�?��W�7�
�!JD��v��.�D--�V��	�b�a),��FP�l�Ƈ1V,�w���*0�Q"�$0��G��ۊ�.dSM��`������P�U�68��9�Q�7) �W9d��Ky#���{���?|�	�~���{��W��a#��?�]��/��T�����쀒�Q�8+}�#��j�`�<L�ro�Q��@ '
Oĉn,:ɍ��SH�F�h�w%aѤlѧc=[u��ϐ�Ĳ�e�Ze?�u�A|5٘m���`e���G�g� B(�t(��[N��ʀ����y���gfc,���I2(�������θI�"��QG� �eq�~�JȂ���P��1�9qh��߰��`�nxˮ�w-�(��#h��wwg�$A?}A+W�q��B�M��A��Wih��m�6��Z-���ԛH��T�}#�=3Y�$q�a[ͨ��q�R����R�-�ϗ�`d9� @?�^�hkJ%`:�X"���z?���l���)Ò��x�7<������R}���Y,�TB�Q3�����A�wwe�=������ʁ1<�Z8|�:+R�%4T�����6=H?��g�*��b����ZJru 8v���Ǎ������A� ��g�M!s<f̵ߚ����g�K�f���b���i�,�
;vZғ5�*C
�`}�<k���k�{�ب�^ ����\$�6�Û# �Ѵf��!�l�2�F�л�q�Y!�\��$���V(�p��yі&�Y!����,H��-(���M p%3����٣?��Hz�C���ʰQf�����ϫ�SvM��D��33c�ڹQ�LǦLX�@��������8U�W<4��4H��֏P�b�m%~�C��Sѷ=��B$�y3���/�R�yf�>�w:n�Xh����(B���A�@Q��YX� ��M������3�b��y��>&�ڸa�GG�Ŧ�����P��X��e6	�o��w�"�g�H�Ȗ\-���伎�g��,�ݿF ��7�D�7E!�F��/�?��@*�HO㑑+Dk��)�_�gt@N�qЋ<=e�	]ؓi��k`nux{�7��z��,��F�����yX�@\� ��R�l�G�Dt
���z4F���y$��Cm(_Aዳ��J�O���Q� �2|A�͟�H}?��V�ax0���TX���Ѿ"�I3zP��oف�z�a=b�_������&�>W��:ү:r��s����"���	�E%]qgn^��ד�3��[S	� ^�d���7�����!�1�a�qo&�Jw������X�j�>ߎK�>>j�/�^5��:M6K���1����`��vN����{�LiQ�+�NaI{R�����":ڌ"����I�x�2}��{L0^������@S�W���3ڸ jy�w����n�������w'ӻ�6f�;�<��\f�g^z����v2ʖ�QT��>�X��v/C�����L������I�U��y)�E�Ǌ	����_��^���`^ ܁w`T�~?+6Z��ȚNM�QZND\ک	�"m�Sh�4����c��+��
ا�D��F��]�����UW���;h�g���^Zߐ�5�IͻH#�̻��x���~WJU��hU����*a�O1�%ʊHW�>�I��aͩ�� ܙ>9�1�9����]��K�F�⚗�K���'-2�Nb�(J����?�������~U�2F2Ԁ�X\� �r-�~-�j5�[����C�_�U��y�B�c�#Ţ��ќC.�ܣ!�]�n>��b�}4��>����)����K+l8m�M(�=������=�;�^�	��^�(F�Ð���5��muˑ�ٱ�#t�S��������۲|6^���{�8�(+ڀm��[�Kf���I�f��L��Ĩu�7���?�?k��-V<�)8y%�Hӣ��:�}�,��}$��N�+p�̚�w�1)�Gnr|����(9�(p��T��g�;�%�	���u�8~�5Bfc�¨��:*
=s�$���g�TW���C10�K<>7�O&���I��/�z�#�- ��v�`.��x�8�%^��-��Ğ�fR���F�V`D��p�0��f:�[�8+�Tі�,z�ٍ�gT�xV��4Ÿe�-#=]S��s&���6[��4�����o�	ڞ��{���+�&"�[9�Y9��B�v��l������8��I������߆MxzӲ�~�����U(�6ma���}:b�Y��|����E�:]����/�~6�U��Y�6K�z,�ӟ�/��Ԋ,sˊ�9|iWw�j�1����=����g�F�ׁ^y�F�V ����J��tb�8��)%T��J*;b�.�j+��}lp48Na}�Uل{��#��o2��%����lȽk�]{���!���u{b+��J{�<>c�;��`�r�Je���>��V�c2�'+*�Z�O��f��HE�%jp��kF�-���6�ͩ-9�as�w�8�g��V���T^�NYG�Sa���iMo���F��_DC5�ER��YhF�S|������t�?z�(����ξ<n�Qz^]�����t���[C��G��, k[���re�,,����"���Fs��Ж�(���#�s_|B���z�5�K������0���@򪝧/)Cx�p�<wj��g�Ҟ��4�H����������|�ї��������*'� JL�E����)����O�v������a���=�����Ho�Q��1fI#�g���Wf?��?k�SB��sv.�U�0Κn�u�����A��g�କ�W��µ�+'|j��
:�� /�{�*Լ�1�e�j�_�o~~(��X/��{֒E}���	��miWpC�ʓl�\<R���d�n]xa抛?�D��/V㋄Â�t�M�X��-��D���8�-:�l3�/�݋�ϖ��u�N����v���e��EB��ySa�y(f�^ޞ�@z���{wO�zȼ.���wŶ]D�D��2�$~�)�?K�gZ;$�\��� ��/���˟_���;K�;'�s���,���
|3�)��]68��<��d�7��[��?S�u��,���ʷ��z��&~�B�'o�@�~�p��h��[�rZ�eaCj���>�>D3r@���	v�q��6o	JCDӽ�FG�S��:��-(�l9ai����A��2�+�Q������]0��ţA�A�:��唙� 0�@�ϼ3��1Ơ���VP��g�R"](\��$DIfMk��L}j���$p��2�σ��i��`w��w��}SĬ��:2}��3F�0X�}5 l�(����D�<�X�~~6�l	]���Iβ4��t5y�"4���%��NE������Iԕ�=/ؼ�������X�����u�Ñba�~�#�a��X�~|)K�G�W��+JBc��s�����J�f�{=(�����͑�� *q��!w���.â��\ZY��+mG���=V��}Cu�����o�G"!��RS����2�U��-����F����[�N�w�J����U��$!	oo�d�����kiBu�UƷ�0m��-�>�Bl�I��<_ʅ_O5ͽ-Q�[we��xW~��^�7=�N$�w�|�6̼�!(�U��Li-�r��J8��|T�M de��g�|l�_��N���^cfI��b��,v�a�\o��b���W��7B�-ZM�#��_5��Ӄ��?�R�aI3����/,�lb��:�N<p����"��
���Nĸ''�Rh�'o.��,s����&b���3Ҡ�E��G�������8���7�}���qv��q��Z����k���Tْ_v�B��<,��p>c@���3�̰)B�U΃`�"u�M���e�����N������ng	X�`r��R�
z�8��c��[��	W��,�7��{�o4���&����4�g��8���p�B�<�������YO@(5��7I9�-��\���j^���3� e�'*C,��3vX1���8` �U�8�)t��g��1�T���(��L�1^8����8�k͏^}^=��_�Z�6H��u�	oh���<�J�%��`˫>�����8,������޺�4:�#�x6�b��P�� ��t�}�}I���6��N,(�O?�Qx�Y�ힳl*�d��4��d�t;�J���{\����O��G�'ܺ��\9n鳦w���E؁wo��^�B^^ދ��u�ՇO�����.�i-�B/	5ԤGS�`eS7;_����^Y`h���c���v��)�t,�WGg5G	�o(+�Nt	����q`nC�_�L�Wf_��қSPM Rh�?b}1`�s8shA��2�G���3�f����j?!��Wmw�Ig �O:��b'7:m��"�Y�o]�hS��a;���x��*�j� @@��6P��}7�jn�4w�zv���H3��	���I�YcG�vuT0j���k��e/L��1���i����J�`�� ;����C�k^�݋C����|OX��uhvI����L3V����p��5���	�xل(r���]m��u��N���5�>H\�}��҇��+x']�U7��N��!K�;��3�v�4�\:�_E��|��]�B���2s?.6�!�� G���^��F���cg���.m��e�3���i����"}�T�Dm0�BȜ��mV�<V���cE���KTO;?'N ����+0�
�3��?Q� /.մT%&�R�V�ӴJ���J%�//���xǻ��WQ7R-񣇛1@��5�N.d��e-�ٹ���N����m.��{X�|�G�%L��N"P��VR�{�}�̠v�Ȃ|i�c��J�ܹ�m�I���w�2,9��*���Ih��(��������������N��h�D����M�[tU4<T����/:!6�-�'�Xٌ���j�~`RW\ɾ�.�{4i�󔀫 �԰V�gI����0�A��*�7�$We�z�Ǒ/JWNG�'T����a顋�uY���ؕq���"x���_Ϟ�gy_�nsTK;��/t�J݊�ĥ,Ol��P��9�����h��Td��v��SIG��u�^��,G%(lE��*'D_��Zr�~f:E��H3�<m���ٝEԅ&'�B��lD��i<)񔖞�z)�N>O
���'�~�����n���:�}��@l^a��yYFo-""	~a�[W�<2//p�|b�����l2i���Qo�sڙXj#dXN�J���3��w�DP�@kLA~���!o+[�3�$�LV40��'R_Wx 􉋿 5r��B#�����g�g13J�K600Z(���Y�6�	MSS��r�%%�T�"aN��R4zG`cf@�W��ٲ�n�2����X�+�ë��To���M���5*6.	�m�{ۦo%�;��m���@���Z#���	��!9N�ܟ?�fB��';q63�~��=�y��o. ���H q��;�x�&݆h�b:���q�۴��������U��d�XO�d�jB�dy�TW������!�]姺s���X��-�\�ᢌn8��s�(�3e���;�=&'�M��6,^�����Ĉ4m(~�(��S���h3����O}B���Vطy9?�8{���zd��������̝�iW����#������D�{9'�d��_ִ?����>�=V&��M���0���j�:����t��͂��~�ÙɅ��W_*R���VY�<Ϻ�gj[�z���K�L��������^L�<����M��Za*V�	,=<V�������G73/����u������Y�<O ���
,7��_pCa�,C4=����[�S/�����R�b6�����k��e����59ф[�.B~��mnn��(�N�Vh�K�Z+��k�͟�7�<��(���A�t����?o�b��2�t�u��S���F���A����F6����QyS"4��
��Z���C����,�%�yt��p��l�l̆�߀��Gm?�L�|��\�~�Y}}/����awW<�"��n�x���~"��҄u����*��.��}�vۜ�a ~��;����Ca����T/�A+;���	Eg�R��df*՞|�m�mu]~��AC
+Y\?ti2��{�ґ��k�.b
Mհ����Qccu5Ь�k��aً���1I���ٍ�p1?�����OpIh�'l�l]�uv��"�#��E���$���v��tX�q��b%DV~�y c;�Q�2��`$$,��kBj�]��:�U)���uvی�z�3)�_]�\�X���ţsVw�~=7�au����Iu~1k��i7Ǥ?@t�mm\D�6�2"��u+�����H�����f�Ӈ����ޞ��ֲ�o{7p��{{T:�M��s��A�'3Y��EB�Ϳ1g�vki��f�G�)�Oz_q�S��fڐ�4?��Mb����o!è�����=hDn�.����"~����y����l�����|���hf��L�#��>��:�TZL.Bo���r���l�'�k��hMݼb�����M ��@˵�s���}�%D�} �Y��}� �'��CV4N�-��آ0*�إ/z��(��4�GyE@|�������d[��84%6���..�'%�p��G�����^PW ٞ�w�(l���1�r��յp�I�S5��►zP/�TK;b>�+��ֆ?�ѿ?���!�݆�T�ʂ�PLU����=��c�M�0C�Y�����E�K{ 6��j�^V���|�̞��,��(�gY���G����d����OH{1}uagv8|���M2��(5i2Ƀ֝I����'��/++Q}���Z�cdl*�"�KQv}ÅS�5T�SH�*$\_׷�bh�\�96�\�oD�Bü�;�\M-G�� )¶���D",��pߍU����քa�$d��E+j(��٫������Ķ �C~��?^휀���������|��9p����6�����Hx�����a먩hD0}:�� 9�����J����N�z�'u��˷󝦯ޤ?�[|��a�U�5NA����G�*�:A��F�����B[��J�u��ȸ+��։���\�9b����xQK#jK1��Sy��L
�C[+? 1Sͅ�[�v窣�YWMBp�m<���Ш�X���-��W
�O�zO�@�猂>\�se����\V�.� ʿS?��q�ع�o�	�
0��yU} 7�5syIiK=DrH�Z[-!6U�x$Ο�����;��/�� ��I����Jb�`%��[ל{�Z�Y�\���`q�PO]8�ѝxI�����2�OB��~в�JCbe"J�J��=tG��2$��w?���F�J��c�q�������/���B��8!@��VAD��T,P�O�@�z_-��$j�N�����*��5������.��}y�^�������*-�Pz%ӥ%�~�:�n�^�! y�Sr�M��t}��Y��������� Z���Y��.�	W��V��Q���u��i�͒Er;����u����U}��42��1BI�Z���(�ߞ�SFo$��}���yy~�W=]�ˡ��j�U���*���t�KHHHɉ5����=�c�fU���iSnf���ǫ��@%O��u��ΰx5c=���Ƅ}�^'>�]���kC�8��sZ�R�l���ڕ���(`
rwj�Z��!6bc�M��~����dG4PLg����3���؝�v�	8u�4[s �����ʹ��TT�%$Bs6���[{�
"Ge�\,ij�sk��R70��Q��
����R%.%���N��㐫&��$�oK�����eC5�7��O17q��x`�y�ҝ��W��I�Q�d�$	��Mt���_�� �uZY[t[	1�9�y�^��r����N,�e�ن��	E?|ۯ������E�{e��a�+8�#]�W����Ɨ�?�^�3�)���h�i�ߔ�����bE��]�R����b��1IA�M5��S]3��c���6�咽��#�E���mm�(xg���a�a�U	��9
�\r�3��ޖ�����8)#�mwPx)2����Ԙ�5�U���Q�%͕�@4٪��������|^���įx��܊'��*U�|d���A¨��/� �-}�z��n����U�}R�݂<'��o�>�t�f��5̽�����[��|i���*�n@�Òb��F�̾ѽapyDQ�����̇�}2P�Z���N3�红6r3�vқOc���l�N�w�d��n��<�}o,�*h�W���Uc�Щ����{�9�ͪ�F��^�<	�&�8L����5z���$��g�8EJ/��x�A���&��y��Ϧ�>Q����"���;�P���1�������a���ȵ�� ˋ����-�.H�v&ShO�[��~����gٲ���&�奁Z�D¾��y�;��0����=7�&����bL3�M�D�g���Ű?��n�Ĥ�a��b�a"5U�@��Ba<��`�����a��0�۷�4l-K6Y�D�`+���B���q�X�Ţ�^/O�A{3I�N����̼�?q-�E@"{�y~���L�l�.לi�>\���*��@����n�_1^�B��M���x�N+/rqVW���N�m���@�و^W a%ԥ"����,�Ʊ|}1;�y��6��ǃ1�x.��ҋ�=t���8��/O3��8�R�����K�|�	��4�e��18jq;Z������7�o�����ev2Ar�ۏ#M3ɩHA�%*�V耰\�;!9�t�ϳ���gqR��2l��|e}r��X���Y	snv��6���r�CVz�E�N|?	rY	3�)CU��	˩���⩉��3��mEa��-zBk�ʰ�9�8�@��i=�Wzq�:焘v �}q�sޓ�K0����pV�����"�B�[����[8i29���h< �,(���zY��9m��w��7%�����wGdƙ���S��U�A�Lxۃ!t�_�����%��/��nv�6��/s�%)u�W�ٓ=�Zp�ºwS�[�M��<��u��e@c{��P�����ڎ}�7$����AjN֩Z�t��0��T���@�����U�$*�t ��e�����D�MNVgH�1^Vd��e�q���!��=Xe%��[��[a��HCy9&��x"sl�ݲ �B�!�%�d�T�*����-@l��Ya����Ů$�.���I�.���S���ol��7;a�E6n���I����1�Lǂm�o�f@���6�$~��h���N�"n4s!�O�$_�
�#ͨ����H%����2�~��@x��7}JE���`����Wm��#e��/�;x��ml��c0�.�CГ|���X	ܺ��'���
y㜉�=ϱ �8��̘B/A�_��'��XT��J�2�&��S\,�B�ۗ����2��&Ò��B_�/��u���{�,���w�ي��C�Swkzi��mw�e)3~�g�e�*�������I�â�3zq	Y�`�q�Ͻ\<�C���_v��X�:N�?tY�ե���`��A�Mǚ6�
���g��x��`LT5N��3���y����=���2<��!�����V�l�d�yʂnЌ��$�U��
��t�H�$uLr*�}�A׮n������d�t[_��� �� �䬭�N^+������i���,.mg��ʨl	|�S�`ȨQA}��R�L����u�z��b�PI�ƞ��D@B�[U�i󉾈m��Nm����t�
'�3SM�n�q��α�xA	Z�x7�ک����'4����+1��1�>��U���`+��1V�����G�����eE\��7?��lt�(d�k��T�IC�fJf��s������2|̋�o�b+,Ԋ2,k�n���O�U1(��VmL[k�l\n~Tb���_�QR��F��5�	����6>啔U�Z�0{-5)���%��Z�c_��y4��/�~;�l�Z���ռz�_Z㢃��ű����L@�a�+Dh��H��@s=Y�o�'�݉��MA6�h#�{��+�4�n�QYٽ�7��P��d��\U�>��Ʋ0�w<|�k��ӱ-��n$J����)$W� ��j�	�
�n>w��\q
޺�k[a6��=�@6�aUM5����� ;/��ץ�j��恨?�Y�o�\���71%��+X�td��<yf)S��Z�2�{�u%;O���e, gRR�-�
M;+P���XcG�ԫ �rq�+	F��g���G�;c��G��Wܩ�6�:����d�1�堖��ҫr��v�A�,�oWV,��J�]	������.���x��/UK-r�|Y	-��D��Kc*J�˾�{���c7�WZ|o`VH��ӾB�m�g����24���H���3�c%m�~Ko�8Mlv���\*�/���\����S����$%�sb�Η�g��W���0���w�ͥIf}����}=�턞J\����1�ԩS����데y/��� �vm\�aR�����vj����aj�Zd�CQW�.��+ ��MW� �����z�tx�&��fit�����/��58��'�r��&�0�t��O9��ϳN�-��痺����j�y�*�8Ŀ.j����Y�U�����ٗ����l�j�e�4��|�hg��.'��G�\����g- �9+{�'m�k
�����9xl]?���Lr~�/�6�̯
�ى�O*�:78���ݤ������M~<y�0�4Tԝ��޻��+X��h,�}�J���!|�Z����n�l8�cLiL�4��7\}��}m�%��*�vl���[��

�����4X�U\�:��E�˜���/�u4��Xߟ����n
��Ϟ���82v��K�{�|uG��������Ō�L� o�7�i�_�~/w]/3φ�����ޏ�|�ľ�v�w\*�gL�ϗ'E�,�q��V�%0��r�Jc"��@-NP���kG�����/8 "�R_n/�/��l��Lî?����{�W�[��/����Ld����J�۬�=Y�6G�x�x]��
��4x�������ʡ��@歵����ز�0�9��N�qcüo��@�]P2<7�7+,S:(IVS<���RӋ֓p�{�H��F���͞�2���呀'1c��@5ak[nm;����g`�Q*�+X�K����tB�~b9�� ���g x�|;x���'��ηI�ڲ���Хl��'��$�|'�,������F].�N7Լ��ɴԮ���=�f�&��G<0`�4�?&ry��_#/p�
�@!��4UTu�7Чէ���1�𸤇3}��Zo�0��{(6߿��"���'��������e�W秛��J=/SI%-]��5?k��W���n��Y�]`�̉��9��y�ˎ ߷g���7C6�R�z�Y��񝇷\��/���)7����%��s�/�:�� I)�GÌ'�Ԡ�dr�a��#B���������n�}�g�ֶ��<y��������?V��_�E��B�����Jg�1�A����7�@z��3��,xt����U�R�p����T�&��Tf��`�>^�y��
�߰^nb4�� )�}Y��H�r��_w�z�&�ecw<�fZ3tV��ٯ���Yti�gS�b��l+�/�f|�ي���x����`+A_N�c�˙��2�O��+ /���ewlQHmB���z!�nn��#odC��a������?�,U]N�K�j�,���)���k�y��<;���28;�R;ɟ_�~)^��h^���h��*5^2�X��^��2��Z���B�N�j���f���'.<���h����F�	M�'��������v��p����A:��ӄ�Β��(}p*�5���$�Ű>���������Q8��ʥߕ�����(�A(��C2
2�f���Z������<����0�����S�(������4����N��r���f�h�^��$�E8���e��)��U�����E�n����R	�\�p��Bn�Q�B��.>�����_�ܱ]�_�k��K�Ψ���k���Fm4���N u̹A�c̱��yg�$� `Q=�+�G#bc�!����]�!	���ԭ���ftU�����qt��/r�V*�1���M�i���:����T5�:-��	�x�-�lFTф�f*����Ϋ�֪rU��&]����TK���̝x�z'Hp�^��t�JÐ�/Y�Qx6��b�W�VR�ۊ�
F׌��i+Lg.<���'`�^xSu�(
����geCa���z��`}y?
�����=MD���>�R�*�G:3k̀�i������-=\㸢�NZ.��+���"��t�^�X���y�p�y}aR��d�]s�>��"��]-rB���DwP��K�S��#B�ys���+Y���4�FU���v:f;QO�,�<��:,���Ձ	G���H���\R� �t�"�.�s��_���爭)w� .��J֯�ʥ*�th�ن?�-+��o��s�9k$0�n��t���+�T����p|�oN�W�ø��#V�0d6���#u{�q��צ��I���$�K{�=^E4�[��͸��Q�'����w�N�! vN]L�(G��jb
+VB���B����O�Dl�/YY�wZ#g?���h|����5��G��Y��n�� �轟sJ1é}.�C���ϻA� �%���bf�]C���I^l)+	�v@��k�����{Ű''�ﮫ�c��딉��Ϧ�UJP�ǻ�o5�Z+���T�����\��I8z#�۠����I����)�_�EFQ:/���Lu?W��Ͻ&yy�T}�c��eVg-\��"DR�j:f>.��;���V�v�������|f�ud��v�o��a~���Fr�������?U�(��6O���#�����g��S�Z� 7���p���ۋjYp��b�TdgBe�gsÊOx��dOk��� 8���eUh[���w��VN��Yk�R�����̴`�JOL8�75�W�L�eT[����и���;$������-���;w���:�������?���v�=׷���m�1ݾ��I��� �t�zoi�梹xs�|Y1����@��x�|-L��ɸ��x���2W���ȯ�xX�*��R�I���]A9��շ޷�jq0F��V�j[���{Vr��[�1v�d�Y��6 �
��:��5�a�QVDA�������������Py��JW����{��Q��>�=6�-��F��阩�c���]��kP�M!�h׭�ʜA�!�����^�S�%��Mx
&�*f�r�4p�d�կFfAS�P�J�S(���p��|Q�gQ��5���F��}~-k�ϫ���E���^ �k̖��A��m��'_�'��7��]��dߓJ��/=v�p�9o�[������h~����e۩u��>ב)�گ��v~Z���~_$����{ӳ�s@��]w����>���+�)���3��?���2�Frd>�y컙zM�2>f��.?1b�����$I�:�����RA��z Qdt�)E�{��Ğ穳}�\r�f*lQ|,kO`�7t�b�;�"�K���h)[6�&vP��̭�HZj��|Ŏ$cIް�~ �U��l"-���q�<\cՁ:~Ю8n�a���W^���z�|l�'�˱�/#�mp����}:#D�k*��l�j�c-"{ &D��.�C���%�'?�����	�:j�Ͼ�:a�L�.fOܱ�|Y|��H��[-�A�|�@Y�i% �W�M ���>+��\{�u/�Mq?hB��4��ؐ��?U�R�b)x#��`�3[Tմ��ؼe�����9��0E�g��n�jq�Nzymkf�ێ1����Nw��e;���f
�SL�T��+Ļ>��X������jSץNL��GA��$�;�w�/'`��i;�&6�����G]����!��k.�^�ٔ_V��yR���~Ua�w{���1����1A�*mF��ǣ�Q���n=!��k������D��Kŗ�����ޯ­��o擼6}Ύ��l���>�*��կ:�T�\�l@�kH���h<Imq�ԡ�7c�Ǿg��e��ja,����Q��>������=�2N�$�������Nx�RR�A��Z;޳�p{��:���l�6���z9{�ǧ��� ��J��	�脸ۏݽ1�/^��U���Hk�NE�V��lZ�ZU���b�s��}"��+|׺m��"�Ҷ�&;������b%e�n!N�?�O�?�(U�w�ٟX��3��y���8t.�)��	�G��"hӓj�Ӟj�N�o+��\[tN��X�<}�>s��ڎ�p�i�п)��_��su�	��obD>]�2Ny4c���l}�a�wR�b�o���-1�+\D���l��S��ZFGh�	�/��#� �b��S6a׸c-tnIdGO�X��k����폿[A�8�M܁*���/;Pը&GHj��ͽ��\3�頬����B�p�'&A�3�K�T/��f�Ƹ����l�!j�N���=�"*�?x)�ٝa���՝�R�+�gbj]�Х�gq݁���KM�eE���Ò���X�2]J� �Bx�K'yi�;rҬ�{h`Ғm���A�U�>M � ��n��GRڌф�խS�u�������a��,�����Gۙc������:�R�"��d�-��E��TL�'�̂wb��m��IOm�!L��x�����9�Qۼ2����,�����L����k�D�kr�z�;k�1��rZ�Bzf�Mx���~Z�Z+���j�/��7_YB�Bw�u�~P+���cߧ�� �����X�!�n[�?j��?�`�lс[�Q�!�ַ��ok)>�/me���2�Ϊ^��[���4�o��(����ǷGI�?��97p��Td�	!7H>j��BO��d�!�	!S�2��������J����:\|K=�1g���chK"���?&�=�}��ɚ�'�2+\nXi֜���ًA
�i*3Not�@yφK�a��>d�nAF���6a�26��紷G��KBv6����;. >]�UpP���Bp���0���ɿ�1&�d�Jhʫ�z#dq���9��|�E5pIyU�Y�8i��k˛a9e=�P��ܰ0�6\�`�ظ��i��m�d5�60Kp�PCK�[��i�ͪ����^=͞���[)j\Q��k>Y1���?�څZ|�g���q��r�U{�)!!݁�<��8@d��,��Q��A�Ҽ�p�#��� ��w�Z�݇>z�Yߙˡj�GKJ&�3Ȓ�`�fV�;�I�jh8�NV,ץ5i{bqͅ$g�*+!�ڜ�XpV��2�+�q�k	+|@d�.�C�?L��[�
��L��5%$��OU�r��:��P��F���Y�ˤ_\�=��w__#:���D:X4���(����tF�OTT�f����#EEYk�IU���ɲ_��Eо��N�γ4����;\��>�y�s�7�ԭTx���:��k>�c~d��D|�̖�[���~����g�%���㻥�ݬ�_��E�|~��zP����o˲�����].3}����q7M�����yD���U�h	=T:��E�L��1��_^_�I��*�q�Ơ V�V�I�)���9��(3i��͝	�����b�Z̅�'\��9���/9�S�������B��<F��lN�{G��̫�藽K�f<��G������"�k
����y\ü��ᄛ�x2�@������ц��|+t�A�D�.z�~[G�b�s��=S3�Д*�k���^�э���c�yL1��e�!'�7�ըm�h���a�߹����¦)���a�y��P���ب��,[��z�-V�otE��!��M���9�����7Vac7p�% C�<o�OA'k��cQ�CH��a�/3�(��e?]R��A�K�m�"߉��G���5���zo$��9�#n���6�J��a����$��-ؘ.8�;o ��sN��&�$n��>�;� U^N��i�;á2��o׻�Y�l�i��e��w.T����xMs��	^�A��U�}R�YŰ*�3Hh���]Ml���?n�E����o��$�齐7��O�[fo�I�@�~�X�\x�@మ��a��@h"~Z�5�c�C�T-�z;����䉸��2�j62>�a�;]m-��Y*����o�k����1�H� N�w�e?���t9��_-�Tƻ?�L5�)>��S�C^h>w�Tw�yw=o;���.ύ�����7�T�����6�}�?�8ݭ��Kiy��/ׯ�<\l�c�ۊ��D�֧����c��p?�Ǿ�ې�5*Me�rYC��=a^u9'F7�"O #�8|9�u��kk�hӇTsn8��D)�Q89L��U��#z\�$�R�g� �F���s��jO��?/���@�i%��6�A:�9=Nm�~u]x���zS|zo8F�[ka�l���������Mp{C��C�㰴��kk���������&����S�~�,��`�������r�$�ڲ�<t��f/��q��s�1�S;j�Ϋ�5I���
:�I��ڕ�}�8��$��p3 x���1%Ԙ���~׃�['�V�����1���9j�O9@b�o������eRRe7��.�A6y@�1+�
���AI��e��D�UWC���sb�q^�������R:���o��l��\�='NJ�>��6}�a�ٹ�z;p������lϢ�G�v)I;�,��*GX�IS�"tH�s˟Y�����.tA�]�o��k䂏)uk�oח�Q��{�ۖQ����AM)�"����Z����@7�S���yK�,�:6�~���N�ن�*Xڥą��q"/0�,K�����Y���K�T�*���޾���/��#����9��# �;<� �cOzj��8�q�e�, ��D--�f��ާ$��>��x��s�[��j��,���Z?+u��������UeU�睎|K<Z��^&/���"#�i���n1���Ԏ������"�Kg]�L��;i���~��L��:_d�l���'e՛;�]�k�Q�*\�l@ӱ��ߦ�����2|���|%�ґ�(�yHb3:���pF��0��1d���XZ����+�cC���4.���-�~87 ���)�=�Dڇ�yr�Tp\�_��@�5^B�)��h����*�W�n������Q���H�Ѐ�U�����r)#�N��B�� ;mV�ff}7��X��ǌd���7�C��D���N�a���3
��TS�6�T�-�xE�����-������?%M��W�}n�����q�?��{�É�]���w$�aSH�����i�6l���H=����u��|{.��/�U֚�T������ve���7��F`��e�Ѿf��ǎx��%�n��L)�H�f3x�*��M(�Q{��0P�=͎ۂ0��=5�r4������ܾD��7�]{�u��#�+����H���n6Ჲ��ETq}�����Φ�dvlTB��qN"���	vS�ۇ}�k
���}�>����i���ȸ u}y� ��4����u��⛢��̢�*1�]\B�p"3�5,�ϴ���,+�������r��u��Z�nń R��\Ѵ��Iބ�Ĉ�"w�pu�l���1��{�/u��-�P�C���R�$|(�3�7H�B�(m��Ą�1d��񙬕����/�/���ti��ȄzPVq�Ӟk�f�2�ڱ#��kF���ta�sV:�V�	��9"�Z=Fh;d�c�89-��7���M��R�xv\wO�+�������!�Z��c�-_���������+��d�m���<8��u��j��������U�̦�����y�2DR��Vt�����m�I�&[P�?�t�z*Hg㝊��Jk<��T�ԍ��p�#�����`���zO�n�);6o�[� s9O�9�g#YHXF@�U��k�}����K��M�P�\x�̪�ӏ���������^4���O�L�3I۵@c?��:/ "MQ��eiSh��q�b3��r�yˊ�EC$�|��Zy36E��-Y��Q�0���z W���&k��?˖����ɸ���O}<|�Y� �?U�ݘ�xb���P,���
�0�!RT�tzlB��~O�2z\F\�sT�����(.OlD��Q�V�¹���n�=i����Y�D����܁�t��t���$��Sv�z����I�Jm�U\@��Ǡa��rzl�@SZ}Au	1�c3ԇ�A�Y��8���Q@�Di�4Z sN��2��U��Q��dB�gƲ�i��nEI���U�1e!C�]�$Ń��IM�͢���!�)����5�����*�QƐ��s<_�qn�u�2��^���4T���AF�O&�s��e,SkJ 3��6˻M�Y�ǽ���iq�������W�T_�?n�Mr�-\Xo�}bq�+1XJ�$9oX�2!5/�(ɥ��s=l�x��)LE;��.�p�Ͻ�z��,��V�Y�}�o��G0�B;����_7�`�-9�ʍ�^�m��m8��6�c�3Cȕ.[i?�-	�d�R!����� �XX���� �2{ㅮ��m��K�sAy�[��NUv�u?�	��t��[x#�-���Ru�ED=H�+�tOR$	zf�Ѭ�(6��ͽ�!͖�����J�Ё��E��%<m�"TS�:i�K;{f��kEA}\7or%e!K��K��``�F����R�̮?Eߟ����L��<��p,�^��̹|�S�bR�`��ʷأ㩦�_�>�l؋�����t�q�v\JC��4�Jr�)��v^�9W�k*��ܻ@�n�C��^I��3�:!qbt05.Lgx�h�GO�3{��qT�3b��$��iq��Ip"6\�PFW���W��b%���2�eX��3�Wx�9J�B>؜^��S3<˔�L'�WO�IFh��e>d3���D�|X `g��;'�J��U:عa��] h�>�����9+T 0��TurZ��0F���	<*Z��20&�+H����2�T�H8�'���+�@���h���ZW3���[7���S���
����@o:��Ӯ�zoy$�B��-<j�~�<VH�1O87>�����u��u�����+>e�z��DJ�_�$Pi����3�ϸ]�^[O)�^LU�L1��W���=��(�b����$�B��s`��^%��<���R�C�b.�{���@���!������/�z�	�<ڮ�"�t��[t3�SZ[�!EU����-%c戏��=���ql�6�=p��M9/{�
��G��Gp������e�H�.����g4�f��͘&T��z0���&�ZҜ��78a����0c�u3�Y3[AQD(�����M|3�RP�^Eiz�%(e�����ڈ^�W��n��u�m	�8&��ڪ���R�榛�@vhH�yi��(��KCW�3g+.s�qJ�V1]��t�PD XX%㓂�e��'@Q��#'I�,������]�I�&���'Ƨ�:�~���=�2��1�5���Z	��<>�����`r�)2m@j��}Z�|'S�ٓ�J��իi͒D�5:�z�ݚ貭���{),fݼ�]ҍ���/��kf�	$��&G���2����΃��K?���_��Ċ�¨������)��s�ܖ���յ�jp,�j\!��)"Y��*?�q�����`�7Y"�����k:�M�}�Է���y56G_yt����씻��U��������}z�ۿ�ߌ�V�a�j��B']5�3n�m� ������� �*H[��������)�:-³�^�}K�\\e��1�T�1[V������ٰ.�n����vY5�ޱ�Ղ@�&�8����M!��?�����0'�ʴaz��y�{L�%��C�FER��T
{�h��/^D�ߏ@9o�!*h��iHM0¿D��<��]��f�R���Mq̬�F�q��z2g�,'��n�W�������͞l~ʴ���ꗮ"L{99��ʆ�x2]���f˧a,I����]�mW�ͤZ��4�����4��x��Z��Jo@��^I*7�����3t&���<�9�;����&�ytaak؅�*�9e.'a��`�w��w@�˃Pn\�P�P��?��xa)E� q�����J�|�C�p�,��|���k�{�]�h$�mS��V�=��׌���e"	�g�iq,�Qow�'v�#S�����	*���U�S<r��5�|�8�*��T�sus��&�ʨB��ʦ�(��XT�������Nx�z�Y J�ڶ��nh���>Ota�jZ=���� �Eb�J�e�����z���nu���m#n}**dM�0�?El�2&x�\����:m��G�Y$ۊ�w1Y�Ss Nq������%^{��>�f�@���:3�^�f�ճ��;=(:h�\J�!6��[��%y�Gq��y�y��H'�X���t�'��ׅ^͑l�������+lh�gƬVƙ��G�� �%�
�����z[-�w��{?��f��)י�&w�(<����|��/�������,��!�=�����6��0�������kw��1��A�>�L�WVq4_��F��ΜS�Nў8��5�d� #ۢb��K_P��&����,�c�r��s���(��`�b��i��i &D��7egmf�IU9�|���ƒv=@��q���9��!G�K��텂��e��?3^���u��~�uhy�w�]���:Gs�IA!%s�2����p��2��kx��U�C�9�ٽ�Yu8`���KG�Q/�����4L�b2)�^A���8�b��B���7���ݎy"�{�3b��&O@0�	��R��=���D���|s�*~��mG��Um�1���nn���@��Eg	������]-{4�#м�ˋ}}X=�+�Љ��i \O��~@$����a��e��cN�·1�� �%���2�3y)8������3�K���;�H��l�'Y�WS�%��ds�j@��܇�������^�hmN`Z�il;(ͷ�*Dg;���(v.$������Jlq��!����*��� �8��&I�h\� J�Go���k�%�S��X�����lԖ����=z}��
�^��4^�L�U��kp��&vzm�l�Xz\�I���tQ*=6�<n&y�h�B|��sr��bKif ywp�0��F��Z��j���:l��Y���J��>�L�9����� 	�Y��9�?���-*VخݭCx!/�����O�D]�Z+�O��Ffr�����寢�o��]���I��fi����v[�jk�]D�H�,L���X�D�YLl��_��P��-�<��Z>QcE��ލ�]:�"*�D�V�2=�ҟ��5J�ϗ���g��L/��'i��5�"��H)Ke"�1�ʇf����?��u	���-m]�iJ0|�H^���[Q��O����vD�-UGurT!@����gz佧&?_IX8��mlg@�������|��DY�]��A�q�ό���9�u�+�7�Q�r@��~}_f0�7LG�!��o+l�MѶ@+�ڠ���'	�y�bv�����%>V����gF=�%=�^ۇ�h1������U����#}�A�8&�E
7?���mQ�F���iɨj��X�Y�;�mf�~��J_MV�I�e��:��\gҟ����`��C���w��rT�
8�~�N�o��X�$�~�<����¶hN̰5t�{��u�s�^�'7�/��!�ڏF���A�����	"{�ޮB�����O��
��b��}�n��71����`�l��;TZ�7��+�=ކ)��Ud�����w�y5%L�M&h���>`��G]�z��ǰ��龜@���(ڐ��&��w�[�*%��7�r¤���t���m����p���M-Xbv|��O�j�-���[�a�f�w6s�����'޸g�ZȐ,kK�θП���'�U�,����𛹮n��	~��4���Oë�4x�x�Vp
�='EU!&�����c�dfn�X�@��m$��L��4��\\�|��=�x���L�9��Y�Wb�W�-�y�L)��縩���d���"¿��a�-�;۬@�/�v�3qS�@��b?֐��]���"(/���m#9Aw\_0�aAB�")B|1@	)`a3|�EPt �u4��g�#q�\c���f�!�1�b��x�����;�P��W :߂�g�ay��0������EK*�3W�A�ߊ�iV�̰�ƫ%��=TN������
'q�h��F�8�GA�JQ4t���>�]~�2x\���v��n�L��<ֲ)\����[t �s�/���u����
c�gG4��Rާ ��7-� ��L(7��7nR.��n�-��m�c�����t3�1�0�^�G�e�~��������Ix#q��w�TǹIk٩�.��wq#�q���d z�֡
�Ad�kO�k����Uh�+�{[�� ��@�\�����2�hm��x�P�v��0�h�.d;j�9\Xj�{�1�n�%$B������6��B0�֟��N�F[�RyJ����.���P���bN��k���&~��'rs)OZ��	�\B����!L�6;��Ez���7�(A�0j؉'c�	P������F�$�����~�c�����2�*4�V������HX2�dɀ'����x�!��6S����'��W~�l�(�x@���hr9��	-�_�	L�Q9I*lG$��İ�A�燀��Q��D]ġ��w.��Q9H�Fɚtc�|�	����?�����c���#��8�X���C����D�Y*1����B��9��g� �m�+�}�n��[;�s`ƭ���M�r%1�m�L8��-n��r�����[u��]6N�����яqX5vV?�]`Xz�&E��/t�3��*i
Ыv�����8q,s���\�S���Q;Sw3��rYpNR9�L�
]�����?*S*��A�9kE�_�j�=ń�����VE��b<�����@nm�h�st�k�ߩ�5�3NKn~A�����hFƒP�
cվy�hNV�c�\`��܃`i}�� ����ˡV��g����fJ��Vt)��	��w��0�k�E'�3\��;)���[A!��	kA;A�����'d���8mI&��p��tt�8��q������'�1Iy����E�f`�����>�$�KM�������qH<��/a��S�I0#9�N^�X,&'�����({t�R]����J��D_䢚@��h8��s�3���G�s�̜<Y���c�oΤ�^_3� =��OJ&�������]At�O]�;�
|��|�e�ؾw��<HmF5����W�[�Fd`����.$�ՠL��g�w{�)���m�~��f9�u���ז�݀��f`D�������h���Ƕ��}?�*&���=���)�k�ę&Y�K��jҩEi��23��v2��/b�<�'����61"�����K���lA�!����L��n������K���:�x;p�iU2sRfBh����p�^��)I穢f�=�-�gz�b�>v���{�l��Z�c:��s�g�k��Pq�(:�[	ǟ'�ڷ�w�s��^��i���"��~I���d���P�"���&�΀�k�g}�9� ��Ku`iF3Bl��sm�����N����XQ6��&Uᔞt�����s�8�V�)����	/�� !t��غ�Ѩ2�f�
;-���L��+�G�jk�2@sX�Tu��b�^�l<h7��_L��R)�:��p\!����閭ߜ��h+J����/�g�}���T�Ie�O��N����D�}+�"�rSF1OT��*�Y�{m �$|t��Z�+q�I!'�)^66�8�h	;ؖ	�L`8�"H� ��������j�����z@�9��wp�-��2�+^��	�ن+�l"�նƼ�+j�t�=��f׬`im"���l���ӯ�:B; �y?�%��,�Vo�.���I��28�n��M �y4���7J��JCL4d�G[���,��qm�UXՠq>̃X��E�g�Z�jbR�2�S=�+0�d�f�x��ޣ���>TȤ�<�X�gDש��Z+8vI�=j��	{��j�Z~�����>FE;�d���"̇9O���)^�ݑU�n[A��Po��ԗ��W�o����Կ8��C�'�9"��Uw?�m%З"�z�{X�H���/�=�mkARE��Jއv?���Y����u2v2�=g���}[��̉tv)Ɇ�4���աa(wf�O�"�� ���
O*�U�VQÊ��+���S�)����RzN�7�M��Vf��Z�?�i��_\�H���Ea�r-i�RP��!l�ܘ������y��\i��ap��?؋����1��!�~�*�a�4���~�bJ�K=��#��ZˉV��wD@������*s�{b�"�@�/#�x:-u	� �P;�*l cn_`�$�]#��D"�	@�Q6@2®FP���[���|#nx�?��ʜ�3�dr�kyA� �����Q
\v�����S��Rm]��{+t)�5)�6�l���(TsA�E��9��G��ؘ������������h���	Zf�YfT��˪8��:G|�+��0��Wu(�jL٘��**����~��?�"0!�'�Oo����F3���_��3����l'� �d��#B5�"���DB"�P/t�̰�Ř��H������Ź7��\>��ւ�~B`�IYҙNϋ����N�����LT�����`������7��%iS蠆��Az�S��M������1\Td�����xpG]���k�2x�h�/U��ݞ��z���*��[%b�}�xQz��_�$����g�A�b��Y��0@��L��!TY!-p�w�YEm�e�)����0��)õ���1���f��Ǝ�H�y~s-�v�T~w)�:wt�Х���#��g��1f:j���.�q��**SDJ������M����T�:�/��"h�j�N�4a��z�7�ܦ�ʷ,GS��"���p'|v�A�	��u�|��Y�0�w3��g��="���̃~XF��y�)�w>����P�Ɉ�kjk6�!�x��R�.����'���B�:�x��V��Ut��C���!�*�]�:$��7�s�y���|Aw+zH���?-'��B���(M�J�E�ߡ�P�1�#�-4\�h�!����u�Q�c��B�S �!^�4Fn��Vn����o�v�G�?PS�ӽ;�n�������s���}oF�;�H����s;Ɋ��n���g��a�<��F;-�;���w��y�;�����W�q��%��aAT���L��DZOA�b��	J'r�������E�h��`�秳�
^Л�O)��̐+�A(QQ����r�Aݯ����O�������·P�ҷ�����IQ^	��a�z7�x�m�I�bDS���6,�G[{�!4n�������Lm�7��u���%�����!j2]��,�Td���w&��^3h�͸�������/]੔�Gl��(�c��f�뗕��CY7��T�&�V�����9~4��_}V�n�u��[�g�W������G�X!|}@�%�4�n���I�D���H�tQV>����:`�&��e�]�W�\p0��8�Z}��0�w���MY�+Q�E� #|�����i^�\�F#����Z8P��^h֒1yn�J*�+�X��8e�o\s9�"��x��| 2sbã�W祲�?k�w.�]s�?�U*���S��K����-�K�����q�U�Q������.�0�y�ɘ]Z�*Z,Yi��.�{ПS�d�z8 *)��r�N��k�a���d���+���,�Gn1o��#�p��&�X���[�&���2�����!%b�#;G��R63%�WP�{����R��B�Su�h���&�,'@�b��3��I%w��A�y>�x�ؘ�gÁ�v�6&{Zk6I�W@!����xGƢ/�"1�2oц	��,���<�� ;N��� �8�����i�����s���b���N���_��>>-�}%n�\��5,��{���7KC��@C�pm�ӊ:��	�i���MhG�.�&Z��X
�B�/�=�Y����o�=�)Z�a���:��Ϩ���x�w�p��e>���'��+<�����Ȇ^�j��;<�X!1�W_�)�#=���Jpq�Z���4����B��"�ӥ��^��ܳ��2X,�=�ֳqd2ۂ�ѯ���Lj��M����j��G���I�/�#���8� E��ᒥו�[K|>S����fG9@�h���j�y5��~(H�+ϔڲd��%H��G�׸ہ����)=l�0���g`
�y=�Q>,o�e�e�D��J���v� P��\P��+��!�L���pnI����+2ϯ�`��U�>�a��	;M2�����^��g����	�;o+�}�R�]��p��A���9�]D`yف��|�RE����:�)�r��Ή���s�ʋD��fJ��T��� K��������>�'x�q�����l
���B�S9<�����6��� c��Q�qIo��^���1TQ��>	�U1�jz7Vw�m�Ɠ1��0�)#D?����.�^����RXq}�f_I<D×vK"q��P(MJf�b>I �x(6L�Pz��\�^e��}XE���U���(�N�_ş�h�l�DLw���e;e�w��y�p'VkF���F�������s-d���=��2���59-���)C��JG/I��4y��"s�9ƣm���	J�^��Z8	�.��Sm��?{�i~�֔n>����]w�W5��b�zQ�ۛI�5�� �4t�ZY^%�=U�����W����;�=�&� j�Z�g�Ƚ&s��.;�XV�k��C���q�M�������,w�ʥb1e�'����|A�1FB��SS&9�~e.�z_R3��g�O��a��������-� 6Z�`�����zY3�-9�����ꂤ�� 
˚ȑq�ed�яڍl���5�����\��W�Ӷ����ݕ:�}��K������|yo�H�-�G�-��CDѵ�/a�m���󮐿=�o�:��R���\���R���2�#�n.�۽�������$8�jn�����g�ƣ�L��c��m��d*�� ����9*��㰵)��Somi'%������KI'xc��{b�9���b(�<?�v䧷T��{�p�V�:}��(���p�aj�BuG�ˆ-���h�=�P�_��R�ߜq��9�^c,
�z-���4�n�Ou,V�x^x�,8���ǥ�'��������V2C&��-ItF!�׮�|'"T�����Cd#�@@�t'��ʽ+��1*�%FT�VR�}Ky�ʛ���Zhg�A�*����hd|U����2%���gS�C@1�x�|�ȍ+��c��4�.��P��^!:��R~��n'gp�˖�[G?�ۛ�=�3��W�~~�UA��W�X�.�:��04vZ%��������\~٥?d<��~���ϡ���oh粩l���� `no0��J��	�h��Z���i;@0��s���N���A��V��sC]�Vp��p��/�lξR%���7��3{H�v��Ϲ�U÷0�.�i��`9��ާ}q���l`.������3w!��$�(�~�A���ۛ]2ׯ���M��+i�	9��X���3�A]P���xL�T�q���2�'����Fոs��i1�������)��u��H��9֔��N�^�Tz�?�MR��rh�ц�M]�0�ե;�.���"�`�ޮ�Cs<�L�Ӵ���s��.9�e��3����՝X��Ex�G����B�W@���u�yd��r��6�*�p��|�|p�9�C�4����������G:t�h��}�Z��vR�D�b��z�6_�����|:�T�1��kL]�<Y�3A`��l���T�9�/�6M�7��m*��)/� 2^�W�E'��q����Hc`��e6@1z��)���6�0�+�S��'�{����������k'�c�|�?�;\!��M���K�Qo;��vi�T��$M{�'`���b�a5*vL��9L�-�J�g�b�f�Ԇ���B,�t5N��_&U�q�J�E��x"#�H���O�w񂝨�9&/�_�}� ��!F`a�����:č#�@���	�7v
�bm�ݬ�u��멎v�z6,_�������t�рd������R�}/$��G�ӫ��*�w�� ��htݡ�b�[�-��5gk�l�G4w��|��b���f�9 ��_^����,�N��A��5,@���:?�^HX�ky3�.���J�
�SC�xuP����VbF�� &仟1Bxx����H���T�JL��@�e����C�It��O+f�x�{����^�b�(d"Y�S����%��2�����m'Nۙ�WЛe����(}?�BP��	�������"
��☄�%�og�����A�D�=G��7�Y�� ��|�Kq�9�����7	���b	����.�f�M�;.��O ��Thb�S~g:�FD^��+�m���k�/�F�a ڭ�WA7zG>��Ԣ�I�KC�\?���Ԁޡ����I�q�� ��h�V����;���F�x!Dr{��\x�;̿=�4�aN0����1����5��ݜ�RZ>�YqZ���8�{B����f2�ʮ�ǲ�Ɇkm�(M)�1��pu�7�zLA�M�2}Q��p�Y["w����o�y�`�㉫��D#�cK��\�p#�o �M�=I��{,jl7'^t��W��:od��n=�P�V���A�m�B#�}�!��=�xt�^�z��İd�O���=��)G�$�sS1�~��ߝ�ȣ��okl��)�!�ymA�?���V��zwl2�q&�/S�X�*�� ���s酵C���Bt<'|`@E(���ݨ/o��@��'�T����b�������&�SN���Մ��6%�y3>w�§Џ=\i�sP����	x���/\Bt��$2T
h|����O����7�M���"�37�j�4l@�sO�S4�:Ө!o�*���X*�ޥ{�l�]ZJ�@J8��� �����f��,���#9�G�R���YA��!w�%>��U����r=� ~�U�/���_
#Z�#J"�	�v�xnW�tX�O��r�j��&@y����=0��@�]�?ZH���C�N����>�At|^XcD�y���*�kZF̠O���Gሸe4��y��]6�X9/�����óf��L�;'(��8?���V[�i0�y�/�.f��p<�P�� z[�y����fF�+��C��]^(,��jDҦ���S��҉.�[���H�.�,����a�[�M����o,&���o��iߎm۶�l���N6�mol;�${b�����}/�NM��u�L�}����"�N���}���J��
q��oaĪ\S�j��������f��3�m�v5��D�0kg�E�kt!�V��?�
㗟����j,uB�/�C�s�#�/+��VcUh�T�̎���/J�|W��_�QG�m)5+;~7�����Y�����^�1��|p���@�k����j:���Bߨ���|w[4�s��O����.���k�p7T����}&A��w-M%�]�O�m�*�QkT�|N'��>�?I��ęE��#t�� t�s6\�����$�Eϻ
g3}�+eٯ�g���w�iK�Ed-��2Ζ��b�y�V��<$��c�� �|c��R����󆔋��2����ݦv���s��l����ݺ�F?���uXK�UҌ_����i����z?�O�-ݒ��g*Gcgm�=�;�{O��e�f
[��Ǥ���P�1TF���^�l��b�}���v��U�7�	����ǽ��׏U]c���ZZ0%�x��9_���DJٲ����='��<%F�ߊ� ������A���o�A���� �a,<�t�f�ָ(��e1��u>��串J��dq��r�r�����pJx�>�!x��c�2��D=���3�������ۍ�hR	�k��|�R�{�q��%2�~ȝ�Ć�I�<*�w}�D`��ak�;��z�7ax��&8���[7oH[�q-�#`5�H��Ɠ������}m:�<d�+N@o�&|��IO���ɵ%��,��H>�mq��������k(�@Ƭ�B-�?6��◻t|�H���"щ-`����kMQB�y��� �1��&|�7=l��If.�I��+�I:����ieO��:���n��à��-0�^�e8fu�4� Y���6�x�j�Ր���d�@x��)?'��wm+)|��'�o\�W�xa)���!R����0w+�1g�g�u�Ĺoo�k?؍��B=�4�~u��Y�uV�Ԋ�F�m��� iZ�;6�{�(�¥��7���E�*�_�؊�ZA%���e,�:\�5ꏗ���c�k� ])�G�{���M����'�����P�̐�rm��a$3����~^�y3��+(�䠠N]t`�u��� �6y��dtԂ�Kh�	"���5d�	B�+|�%5�}1!��El��)7����D�F��gx�̊��4���&A>X'��a���t��2n.������}jgXˠo
RK�:�7͗��$�����q��9��������OX��<t�fz!d	ś5[���IT��L�\�-C,{,֑]/�\&:#��"��B���.�BWʷ�<��蕱�#j� zU}F:�9g�j�"+XI�f��m�!�7�2���[����B�;���Ϯ��"CSy����9z�F+Ǐ��S���X���X���w?�O��GPw�+�r�u� ��(��G.Ф�DA5_Į� ~��ԅd*�����5�%���º��7���C�#I8�2�W�鑽U�Ovb�ѨAil�s}-��ܫ?�1x�JR���')���]�L�H�=*����F?��>�@�N�w�.؁h���qkYg���|]&�J0���t],�W���s`���P9Y�L���;�߉4�h_�Wn�M�u8Y�������%�%����+��~y5|iw q�D?�����H!�gD�����Km}���~<�X�z��n�$�������@J|�X�E�����'� Aj2�5�2dÎ��m��2�8�NO�tB�~Ǒ��/,ZI�>⩊� S���3����2Qo��kk�6-����/�jw4�\ 2�3|Q_Y|��@��Pe)����v�BD]��f�T�D�4�Ĩ�84�� ?���r�V@�>.r9���ÜO�9����&S�� B�a�9�*e���w��:��;�w�3|:���� ʹ�Y�s�1��.�ҹ߼��V{L��sscm;5긻�v{Gx=%�ZAJ���oP[R�x���ZT�2��h2T��f��I��0#�� ��������'���ĔM(CJ���^+���q��b� ڏB��E���:��������/>���q�����Q�dQ�,��c����b m[�9����W��{�n�o��"�U,�"H ����a�Aų�(KO�]�v Ǻ-��%ɺ��a����U���r�$�x��L23�
�7~=��^?��I��y��n���A�!�d�����!p��\\�7o@��xX�ܢ������Kε����QVZ���J��`�wd�)x�ZK����>P����ώ�O%ċ�ſ�e�e����;�����z�,�d�`���][͕I.�[���7
y]�~[�ebn����s�Z�[�ǖ�J���o�G���܉�_Oß������/|2 ��谘>����RI��ЙxǮۉ=5�y����'9�:�U2E�;ՒP��E�ǟ�W,�K�Ł�"fۺ9�s�6۔�] ��^	Y~��b w̾[c�W��o�F�2LƜGl��F7�@��rq�Bg ����,M���t˧`+$gyw<���+��N>�7�˵�aŃFq���?��
���E}��l,:s�4E��X��],�iT��v�`=��!X@��cV�iA����<O���'����I�LcHR5��_f�Ȕ�HaD��K l�9H�rI20>����v<����I�WFIwd��g&T�L�:��j�-�H}1�m��Çty���+!,TB9�	h�[��c��H=c�L� �
}F�����rZ'��D�;�Gp�C䢮Y��g ��2+��T~K��m�����6�q�p�xz=@���`R�N��C�ݵ�%t��O��U��W���`��q�c�;��,�vQ׬7��~=KT)D8*�Q0���`U�Xk)d����R?PF�j��n�\�C��Fߟ�Fö �?��j��l�n�����E"�T��1�3$(2�<z�ҷ��}=��wlTe��c NL�/$Y�ӕ��џ�S/��1�,�8���`Wj��tҪA�2��G	,B��i�\����!�K�w!�:Imƙ��[zUڧ�a2�mvፍ����&	��v��ȸ�YF�{~O#�x���m�����m��FƉ�R5�O��Y7��7�|�)o�������e���a��۷:���דH�+Z!j�u�K��+��{g��rYW+ŮL�q��XnK��4dP���N�#k�̫;��/*XgZ]o��X2��u�_&����,�$+�{�u`C�K mU���]�_�!;C�fF���F�aJ���1
�?5�V`$6Au�����^��9����)�Áza+�ڂIxy&�p��lӅY���
��ީv��=���N>���=�ܐ Z?SkɁ��C+K��ꊑ۶�{;6A�f[��nD:��zd�AB��e,�x#�D�Ƿ�����7C����u!H�j�n�^��L�)��Z��q��;�W\G�ͩ���� 3�	V����+�3_�^��*0�����6�<�,�7���.ND.ȮD��������PE򃞎Z��&$�i��@�����X�*ȥ:>v~��\���^������^�Q��һl|
b�ww/"x��fY�YB��{����n�vŦ"o�^d���HH-��T�$���?�BVD[b>�+Ky��t<	 7iA��9�Jۤ	v����/{��@?D�/�%����U�����)�^��-�:�zB�Zz��}�b�2��6��t��UI�6�=���A�����;bᩤn��ȑc����)}��a���^˅�ǹ���>�	"7"{5]G�O*99�/���}_iVi�uD�z��X>��,���C�>J��T*y�{��:WF>)U�'�l���p�����<�M��~���Lr5M���
��>�L�>�r��ybQ�l��u��6D�B�ʀ��*�#=��O)����*-{o���P{@\��!��Z�\�7�o�˾�1��{�Ѐ)�֜o�e0��$�:��#��M����@�;�%��G M`�k��Q�NB�}�l ]�r"p�q�3ő�t�M��SZ�́{�]�ȫ!��_R��)��)\�3�z��sk�FU�c����	H)�����j���F���mX�a�e'��
��zn<=y�w���Έ�����-}��A�{T,��ʕq�Ȋ]�Cm[9���4u�並i�����;����,�g��J�mfЖ���#�0Ta������,�NC�8�c֝��V�́���I���W禍�[���_B'8@� q�ٱ�b1'�^M�O/8 N�E�O���N}�I��Q���'߃ �\_C�Q���)�]��Bu^H�C���b��y���n��Ī����O�l����� �yO�Z
�G�f_� �K��⃏H^,폰�|����H\!�N�Q@ �����Vs1$���i��ߤ�.hM�����DQ��]�8k�d>����L��rw��̃��e��⪚?đ�X�A��;���	Sl-��}���z4� ���^;r���,J�B�/�Y�&�F�VB
��e����]�i�����&�g���%l�"vrs�Sݞ�vd#~�?%��A{,���[B| [���ojΈ�O�FbX��b!��7s�$Vx�	l��N͕��|�*.�OK�5i�W�KJ�e�\%�*���g�+c�eX��zz�n���d�_mǥ�[Q�.[LtwtkBP�*m��@�S�� d�z�Ը�&�rH`�,�R��gl|4�$��r[2T�KHo��'�Ք�-��,ࠏ3yR$�!pxӆ�B���]�e&mM����kߡ:��Ȧu����-��U��6��I`z���yyy���M���7֖(��`=�����p�A��ra��@�_O�]TO59���VDY�� �z���r��Ф1�tZ��Ua�zOk����c�ߛ��GJ�v[��=!�D�*1h��p�����F�����=� ���D����)��
�2k6:���p��_�|������c�hрe�B����lWrծ����n��|Ѹ�p��@�5{������V��H��[ޣmO`�ϜP:0��UW�$o���G����i�0tg~Uo��U��fI7������0����1�0���)IJm0.A��	���[A��ඖ�Ɨ"=����}�����c���X.����Y�H���
f��l�P����(��J��eS�zr��[�g~D��X�����No�|Fb��q�X��Ǌ�28�sRםh���G4�YH���4s�a�6�fɣ$��-mrH/�%������e+�R
,���DR>)�����R[�,a���snUr���T��U���e�egn�9���;S$$�ec��%�s���N�:T,>� ��~Mf�	�������[8	cS��yz���8Z+����*p�f�ش]YH�����ޘ<�o���� ޛB��2��GV�~�/��/!r�e-�?^��́��8������8P	�Hs8�!����2=d2N��7�)��k��vg��S~������,��,�_�C�18:dm�v~&)j��rT3/D3���?�G��ߗ`8`C"���횈���2��µ��x��j�Bh��<��U&d~0Y����Q�4v�n�Qb��|�vY��:>&I����u|�*t�!�:�,���}�Цx7�~�u�yw��\akPux�Y�ͧu!6���� ��ʘ5�S#��x���=>W\x�ۑ����uC�
=<��0w�����֖�'����jk�%�t}i�ٓ�qQ5�f���b�0rr~g%��:����@�>��8�iOΚn��A�><]��u��4���"��(2kAu���<Z\�Tb�9}򷮧:0�	����7<��%��<������J�Ь|XU�����Fr06��!3�U��?��Iy� ��6���9�k�k`�ć���řC�ߋA����;�KJJQ�/�� Gi��kh�Ԯk2�^��^���_�n�n^y�VC����~+������!��ק`���4(���1�C�Hr���鶳�Ė11\�p�'nhvdd�"Ͷ�	6����1�$��9W'V��+o$��d��c\_:fވa=������'��E�3n���);y��Z���>�ڇ&\�u?˶��	��T�l�����9���槟-y�cs~#�݈�d�:\��/}RT'��=}}�M�w��԰�]-5y��a�w�B�>���z��==;����~t�R���������g49�4�(A���,5��d a�r�� �R��4�k#Fv=��~��t� }RX��1�Ġ�# �/�%y'���A~��莢���/���|(�J*p���d"�����q�sۏ�K��R��ɴ|�k�(1	���SLX+&��
M�8�������؇Hj$B���~�yJEW�S��Ќ����%bbn��QI��\J���F���D�kS�4ݪ�TKt�8���>�\|Wd�k�G�"\���+}Y�?Y���E[ߣ�U���@����d�KwL�UL�\�~J��s�l#���Q*\Fڲp���nk�!�Vҁ���ɪc1hi9���j�b3���;d)l����"��V~{/Q�G���D�0���U��������8��m|<O	�6�Ud*a%��K����]L��TK����	�x��m6)���pQ1L�
D�ۖ�:�,<x;Q7R�*L�b  ��Ϟ"�m��f���w6��K��U/�3�������ǝ�,���5"�J�w_��6��Q����W 6�5���!��3���{��֧��fjo�n�;�x��b~5c�F.S�4>�WA��$]�w{�T9���(?��r�X��J]�q�ۮ�8�5]�z����/�o~tq-��鴼��h�Aco�(vvL�'z?K���y ��}�?�>*�L\<\U�70ړ(]�o�'"����3����������d����w���{q�NR\T1���K�������%Έ���z���R�Z�ͷ��rR�:�^�j�W?9�#TRPp�^$^u�l�|�4��E{L6��el������)��H��-���x'���	bs�7�w9
Tm����"@��=N�9����c��R����|��]�e��������3%n8^;G�D�N��H������Ū?J�0�D�l\'Օ�^�����F=;R�t���B��Ɨ�y�����Sp�E��i�X� �� ���7[�J��$��Vs��ѳp�����-nI�{/��U5���6��* ��5��C�,:J�u�yUlu�bȭ��١�� �y�ƀ��v�!�u&��닧�p�4Hw�RL���7=6��V��!���U��B>PM��ԁ���M�{��"���ʕ�b�B�������dG�c�n��M������3[O��?�&>�F�]�%F�k�"jM�\�/�T��l�U���C�#��SB�R�^E���o}(���H5,۞o+�{��������4c�6-�9� +��a�l|vO�C;ly��(��5�W}ҧ�(Z'�6,C�Kw?*K�:�C������Q�p�_m�_-F�"_LE�{�D��A{�@~�߂�6R�
[Ä��E�~]� z�G(��i�fi�������׫х�XN�׬0i~�l�?�FG��T�RRP��N���e�/
���*���7��	�S$������K�fϷ��$�
p1�=�2�tP�㛧����V�"B�'9�8Yn7a��/�-����m�p�|���j�J���"�ו�ݒr=A�7��*_�i����@���Z;�у��G�<Q�츟�F2iQ���o0�f5M��у����{kps;|J�B$z���l����K�����!j4���ƞek m��oc�N�e�ٽۿ���P"��臱?������k�-�)O�9�Ֆ��
��zI���Ĉ�G�5h-]p�ȴP��Ѻĭ�bH�˪*��%hﻗ�7+/�YN��oi�)6MVk�zհդ?.X2��o�p;o��������x�,n~��Y���C:�!X�p�:��P���	0~id'��Z�Jư�#��{4��2`v4łm�ΟQM7�"�Sh��NAI����A��
#Vh-�~�}�G�������C�z�5��E���W�sgZ�{�ǡܳ@ᾝ�܏pSx�z���%���,iP?�'�Ϡ#�G�)AjД�چ��Û$���<'����{�k6�I�h��ا&� ������b�P� ��?b��/��E�į�w��0a1���\fl����C�P�q��>�U0iJ{>U���b�E���	٠n�|����T��E�ڎ�jQ��Κ���سVeb���ۄT�V�v�^�+o8�&���~N}�ޟ3�������ī`�e�!�GӞWjR�RX�]�`bJ�u3l[����S�F�d9��q�%���<��:�zI�6�GG�G�Ю6#3���P��͘�|6��睗�%2Ha�|��&�Jm�$h�xIU+�\7r�[j"��cQ-H-��i��N���B���Q��$�LB����U�:���Z�[�(�vsw���)����s<-�	��OV3��̔�JcR۴��I�#��
�Bm�ľ�* 7�B�}��i�B?���F1���`��2��s���I5S�!��=���~K�F�k�ϡH3-�GW�����e�����C�Hv;?�j��>5!�]�A�]!ӛ:��
?+*�gSծ>�~�~�,�����IV�Lv>n[>��#��QƧ�Up������
D^�a��z?����)��?[����1@=���^���"���S�'�g$Ֆf�MR��v%s�ճ�h�9�URh�U��X��F���4��G���.�������j[�$��{��h��!���׋������~����mv_�U�2ҷ�?:�#���p��f�%z�V��a�ʾ���zӘ)�ZR&�/C���CɅ'�Q4�mh�Tr�f�z�{2�e���9AE~�p�	�&�<�BԠ�h��Bd�ş��п�u(�jl`{�	��/1���u�|�̊���W˯�n`�$4����^JΈc�ӖrI�e5l�g:J�+\��tgɷ����>t����"�B�L��Ӫg��\��4|�p�:w�/��,��_#�{�Dn��nAσ�%��\��ӑ����6�E���Ia�t�p!`��̨��[�^͜ �V8���X�o\!�A�7e�W��Ч�ko�W%*��fJ��g>d[��������U��0�sʆ�$�ܐ�\�}ܸ�ؽ���I��B{$���i6x}c^���k�y�LO|
����>��V�{��fJ%��h���߬����.C�F����"��Ge�	{0mĶ׍�c�qމL3�����ï1e�G�-��P���r�e�B.��7���z$}�,O�����"H*ژ��Jfz_�0J�pQei�n$B�>�N3z�ظi�)�b��~��ƻu ,��'<䜄��ӮWUL�9�FuR�r�H� �c�Q����ާ{�����y�@NIܛF}̞.��sQ�0u�XÛ�Y��
�jY�I���q�B����v8�����|�h��(2P���+�?�-���o:12������³����5��T��=u<�u�N�)4\�}E~%u^d%��J+���R�'.�x{~������Zw}W�����r6���H/:�k0����d�Vp�;������y�͆�K�E�4G��^���g�~
��q
�W�������P����G_R�l��x��@}�5z�|�.���+/^zX�%�,�W���~�	GR]������뛊	n��N��Ur���_�>3<F�Uh��y����|��ʈGG�������-��ӇD�_�IHB��p#p@,���䈖
\
n@@:��Z�Zhw����̤�k�y�{��_��9�n �[Y�{��Au��Ym�|DϺ��>���U���9_���q=Q���%���~1 ��>uM�(���R�uts>��S�o�h���LU}9�ԡ[�.;��t�����p��\5��1�w����<�J�p:,��p1���*�C�ݰ�TH�:�������LJ�8�W�����5x���LeKȴǜ�x�-?9��v#g�Wz�Z;�c���M�մӧ6�<;�Tj�cU�݋���?��3g�]G�L��`_��8u������V�q#���g$=u\n�˕�Dx5�@<� �4A�j{�/�� ��g�b�E贮��W�	����.�7;!���/$� HM�Oa%��F��ⓤ//JEw��m����s6�`a���b
cd&�'�3H�E����[%M�;n-S��1(	qs�q��;�8��N��{*�4 ��_��.e&�\��Jo2�8i�:�	@iB��P)��7�����7#��F=(�x�By����0�L��L�^d�N����r^��BW\���Z-���WBc<��*�B�\�~���=#v�o�
<���k�:�c0�΅H�e]p���	X�D�<)F�$��.y�i�r�q�|k�bh��@gvq��������A�?�.��Kh%�q���GvA��?+���}h��1������|O��w-�0�ꇐXp��`����t�υ4����G���N��[��@���
9:B���A^C��6Ȫy�+��%��:��zO�y'ܠ�f�W3�W�FB��K���&-�o.������|���<�w�֪��!)�������CT��U�!{�� �#�J�D�4l9�{���to�C4]�uCY�8$�|\����{M���0|&0Du�Wr�� ��i@�.��Ψ�'��ޝNO'�5Do����dq�K$Q��x��P)��9h�hi��� ON��H�W�m&��:�0 qʺ|X��+�T��86�6�<#�'h�F�6��7{��f�	�y�Ѿx�"�6��C�L�NL�Veً�]'�tz3{ei�Ws�!B��2J=gk��MY��O��nGbݗY�ڡПx3���xw龜3q&QP{���q��A\b�\����.�eS/�Ѩp��vt�NS�!�c�.1圕��S�q���3�~�������bh��G��ɡi�y�u���#�����dL��O9�����;��	!C������x>Õ#�y���,���S~�_Col���k���H�~=��9b�<�����?���SS+�y�^����С�+�d�|U���X$E`Lݚ'�������Y�̲c6��j�_v��Gt?O:N)P%"��Ε�i���L	�G�"��r�z��P���V���H���[�HJX��gH�c�|}�+�FԳt�L`D�?�	�H��%��x���8�ᔂ��-���[�]M�V4�8
���n��R�Q���('B )/8�f�+F��?r���*����@�z3؍�o�6�eNU�w]�O8Qm�0M��/:!�AH���|Tݩ��@Ѣ���(\*�$����/;��*��p9}��,�dQ��*�Лξ#$d<
"lM���-b���1U?����V��
�3�Mb�!�e���u���m��N/��%էA'}�-��TђzD����
 ��x�5d�:� �nw���}�n��<0�����l��CB��4-���_������@��z�&��XT���E��Z<||����=��aP������yK :�p�� �6ʰL�Ue��=�UD��T��N���:Z_�&j.N���y�W7��̅���/�0���yc4��-�#Ax�?��� ���,נŮ�e��!xķ�7yY�Nш4�(��� E(��5Iz��o�0�se�sG[(�u��Fה8���^Y:����K���]0�)��8��l��6\��B� ���%�<fO��(��4�SЇ=CϼumC����9�����9Ê�0#n]�'�(��l!��d-����3"��G�0#%MA��t���i�7�7$j��M�0҉��e��	�r��;m���᥂O������]�\8�b�~)���V��T�D����TЈ�MMӭc�JõJ���'1�m6��?'��7��S*d?�%5�Q˜�������/fj��w�Y(��t�~a*ә؆:�r��)=�4��܁�X��K��ax�pܱa��^�D����n���G�xXQ(m�?v":>Z����'��{�l�����2���W6ڈ�����@?�(n5��Tǟ��6� Of"�.�x\�d���A��Y�}��YwA���Aӌ�./^Z\n�B�����i+J/�P�B�ņ��d9Re�!;4.�A�3�Bt�mU���չ
y���M��wz �$
�8��9�S�CE�ov���=��],~Jr�	^�^ȣ�EJ��<��e9��`���D�a,	|��a����tn���B1Lq �ٱ7��G+�|���7N	�i��9~�
n+�q?@�0}I�k��D��=��L-��v���vQ�
&�?�ЁH��6�4_�3zx./ʗ�i�>����ٿ;uh���d�G>�MN@R��Z<|'Pp[��*"ްr��h%���=���t֡��ռ;��ڪ���zC1Rz#����t6�̈́y�ó�1�quP��@&�ص�ʄ[|����3h����a��}щ�*��|md�����k���I�on�,�F�2�A��#h������CO.�t�=�hqd .9�R�������tm��ĥ�#4(���I]�c���i��gep�����a@�ͩ�O�v�a� '���/AO?,��t��|��	<~ѽ�k�/�kwB��؍T�?��\�c�?�O��ۖ��U?�L�Q�z c�ݙn$��D0Ɵ�ً���E�D�'B�2��Ȗw��X{6]+1�Ī�,�Հ�ng̐0�#�Ӵ��,�u�JiAF�3��'gm<}�������0'X�c3P����u+���Cn1d�ֳ�?/u��zޠ����_Wh�Wk4��EN��
	2N��\��U�-��B+R�1r��Y٤���=�]�/�z��ơ앥�!D%<7��w��Φ���ɋ�J�y�M���a�K���m�}�����) ��ٽ�Ve5�HSG�5"/`�����6�dcGH�jP���^}���[/p��c4J�;M�K1��a��u���'	Z]���8� ߼Y	�������\G.��yfs�8��kH��ŋ
/����)�I:�A�W]h��B�E1)9.ډ��7�|OP��e�{�H.�7��cn$@��7�=�R?p��W��O  V�D���-b��K��Լ2�j#��x�h�,��kI���qQp�%ȲU�8�Gg�?�z�v��iZyP�W��~�B?�õVʼ�1F���RQ��OT}&;z�j���₈`�����e���\>�r�"w��ǂ�;�����YT]������k߁=U�~h��6����1È�9�%���� �8��^����DW����OA%���r���\l������-v��O$������n�5k��fv�j�y(����v�~N��[��n#ٺ>^��8wY��h�·��̆q��0���Ш��D[�+	�����N��5����)O[��O����}V�L{���X��ы��I�=�+ ��m��N�E+t����4-��d����隗��[T�0n����,�G������������肑�PЋi�m���v���������]��#�T.^J�8�]J-R"�q�Оf�O�����x��^bkwŃA�����"7�&�>!�C���O�� 8��I��;Ơ���u-�r��y(��l�+g�G
8�����:Ft-I�j;2�6o
"F$�6��VN<[wܙ}V��3��Ap���gq�nˢA�HK�<
n^���������E�O3"
<�uc��J�h�/p���c�L(��+ǣ&h��xtn���Ҋ�#�*���W�R�ex,b�/�-?�n������'�~���;��^zb�(��<(��=ݸ�-�"�|yֈ�E�G�9�00�U�[�A��!��֙���EQ�:9A�~�f������`����r�*<&�U�W��8������p>4���_��� ������ke6���+�mG|���2�\��y��3���mx�ް����y�N$m�ۭ�ť�����z����j���7�ޓޟ%��e�I]����|�9@�݂��b��w�溺4�B����������Y�}���Ѳ�j�)c��\k��/%i��i��+��V��O��7�{<W�D��T���$�!���ot�[��_��`X	�A��nNGz��<SX���C��+_�W����	�!��IS���Gx�'�&���'�PF����\efyX�A}�Fn��(�s�}!8~8"��x�9���*vB/ђ�J��*�^Vpa)4�pE�v�8�<�� �"p>A��{26!Ma���6̻�0B!PA"P&V���PѤ�h�RX�^�^��M�w�)��@ٳ�����e���g�0�z9����� ��_�C�㬺N]�I�֨�?�L�5m���Y^T%�|+�Y	� ����?�	t�=H�B�E�7:$Yġ��$�����.e��n0WϏ�`�*�?�t�ޓ����%�F��֯��y��́�dg�\��ՙCluWw���8��Ipnә3�su��`�1��ݠ���R�,P �_��~�i�z�2�&;>���:�*��^�:��?���%E9ɉ����Ӱ�Z���:�����>ٻ�sg6}�ǟ��o������!m�`��2>�<3F���D��&�_U{��`*0��9	�����]]���Z����B�ӚU����MkyXi([�ׁ��ƍ[,k�b��'���A��c��A��A*�>��Mc��8W����.��Ԥ�J�F�[x����j��$ 7���G=��.��.�_|a�^��֞������2�Xu\��tG_����Ҋ�LzŶ�������߄<��h�9�s�jOX)�Nn�a���cb�F�Q�6f��@�U~�%��2��-�㪠s�����y$ ő,l��YW�!)��=�Ѱȉ�w}��X2r�)f11>ķ5�G�̥V" ���쾢.L��X�\~�0�ܪ��ai�)'=�T�z�2^����A'[�t�'A[�(���w�-�-R�Ό��.~�'1�ӻ���ޮ
d�B���я�o�wn}'���v�~�:XwR�vLJ�w-�C:��$?�m{?��y��	H;�h�Z�Q�ѵ1���B�^�qP~3(�&�K��x�.d�ױ z��>�ޣ�m�Ԡ<O�j^?K�ǖ�N$$8;V�D��/7��� ����i�T�D���r�@f��u�+pg�8��[��ډ��w�,dm
�����|�_3���bؖ�ȵf@#��gć��/̅�-�8��'?N��l93X��.�^l�g��\��l9�q���M��cAMPx��k�9aL�H�3qy�1�L�0�fB�@
j��$
r#Z�ſXۊ"��)�߫���,ß!\��T5�b�]��L�JW6�A�b��%=��:o�����4Ϗ����5�s�ĩ�� ��N�d�̘�P�G����(1	>[�"G_�:��n�g �����Ⰹ���KV:{�iŭa!��䠽��w��n�������oX��⌝]�{W�1���d��*�-2���-���+v[۽�����#����F��gX��
��sca;�������x>���/��^oH �+þ��Zc�?���z�σ�s���WW��-�o��c28Cɠ~'NWs5P��-��΄VB�҄��D��]�U%˭_E������{�c�rA�Δ�
�nQj
Ts���Y�"k���#��~za� ����c��&	�t�G�i�<��~�/e�?#��B��k{ZB��A�|��p;a��L����g��6��|a�����r���+��/����T=���q�~a�b���zV�COIjS��x)9�$�P�0��}Z��A*�}����k^.X����%��D�D5�b�#ތ��ft�z�>1s�j�� �v����oih=?t�l�0v�D
����h	+�CYl��/M��c�����J<��T���K<���sЖ�~b�����Y~)߲�}G�?�^����=)
�:�غ�6,�UO19��ͻ�n�P��Pe���pK��A�^�K�[��
���������r0������[Ֆ�.f�ˁ�����c?��H�q!��?F������|9;���S�`ް��9ֲ�8X����8>�\^���'�i󝑪?۾������m�J|�����L�J6���������31���H����+��?ck@�]-~�^���m����x�PA�s����QQ�T]U@Tm����CR�C���������AI��!�i������������O����~��w�fs�г�����b�{:C��c�-OU��edB�4O���˟�}��&r_�����u�x�r���s�|�X�ƪ��aN:FP��:��	�5�1�F�<i_�q�F���@�ր�j
Y=\ȵ&;p߅�5�S��������D]$ @�x�K�j�Tm��#hKOgX�V�Đ\z����������B��?2f�7�B:<Ȭ����Z1��Ey�9Wq��R%~�5D�z����%��y>������V���u5�����2Q/�0_���8�����]�;��+䢏�T�nTt:D��s�R��+1g$�D�g@��������_�T�}��J��{s"�:�Q�b�_�%�ۻ6�����ȼh(K�+�F�v�������O GaY�Q����]+۽+ϖ�|���>�H|n���@�T#�4a�Tb�~q����4��,�sXN��T-���I���1N>D);��he+}(t�����&���Hф/fäC����e�R��UT�;+�+ �no
���4D��Ӎ��^Ž�E���PJ���{7)0~��َ}����K�޵2��K߮���c������O%���D�~��s#xme���v���ݦ@ğ'�X��`��~ι��r��I�={����9���r,()b��=�O��'��s�\D��wn_',r��\�|��2D-*�,{z��R􍋅���������l�����Z2�q��ψ��y�>�J��K�^Au:J46ӵ��ƅ�����~W�"��̓�Y�4~����\��%��7f��ě���W�p1�	�f���I,:�߹&�&8{lс]���LV�F�%�Ł�64ck�����"�{I�DN�����쾉��S�z�|7g)������P
�H.)Y~�$���[	p�*�B�~�]�b��,���<��of&�O''e���Q9��X�o��nX���I��N�ag3�Av��ڂ�HGֆB��K�I+��_t�ٍhqXK�MS���Ԕڨ��R�\J����VKue<��u��~��X��]����Hk��|6 ����O=��l�@a�h���,rjS�������̏�+J�'���+s��>�'p5Y�Ԡ���!O2���`-fo�A�����i����$z��5s=�uC��l��_�菔���r��
����@T����.�){��kw��}~�b沗�Cz01P��Vh�;�姕Iw��"�����~���/�7k�r�ڶ���!=�M|�,��ԍN�չ� �zj�:�K�� 6Ώ��&Pý�4������c{i�z̏���-�ڟc	��J�UF�ABPx�Z��蠠��J�����]@�x�Ͽ��k�SO�E���]�9P�����E����қ�R����N�/Lx���Я���T��@���XީH�UH��w�o�F͊v���
<��'�����a�7�0���$���|-J`9`�r�h��nܽNŹ���[ޗ�n�F���������i&n�����dG���B6]���G���ۭ�����zfШ�L�|~��+�3�=������|���X~�9���9�*w��ߋZ�O��H�W�4�&
z�z�E%W�Z_������m��/��"�+Ut|�p�(���9,i�������s�6cF���� �I����{7��~Q�~�.���dyZ����dw~�U��!t����`
N�������7O9΅����ᖟ�C*
_=e�=6|&*��4���]i��Ɇ��(2�n���;|�I_�3�|���kƊNQ������"j0�h��>�K�
�ta
� kb��xJ��������tr�Љ��;#L��[���a��G#��S�bH?aF�����d�![&��槡r�}���]t9D1(3ΩmZ4�1D�'�?b��&D��9���E�v�z��T	&�7�\�����PI��j�Պ��8�����٫�<u�v�����@H>|�~��r��닲0�9g�����:�Z��"jO��d<���L�F�d��g�%����,Z�[-����IK���,P��d�gn~E�0��W��6��D1f"wDRؗ���I�Qv�K����7����\�\�?a���X�Z�'E�����h��74ߗ����#�v�w�L�M �*������#��b�&�T���m- �� x�C�ۥ��2�I�Ȑ/Ә�������t݀��|������?+\�A���X�S�x�.7=q�B��)"]��:��B�oNB��e���]��q���o������ ��@w���nA�3ԏ¤����O��g�ww��Ƿ�B�w��ύk���&*-�P~J�d�$:�7ܳo��Ϟ��f���=�<Yܴ�a�r�Ğ��"@��z��w^�S�� �1{��?gy�1T����#'�p����r��	����P�zB�ʫ��N�����s&����kqqb$t�ͪOh)�:1��=5��?�����8]*�*ꐔ2����6�ϓ(���՘�l9�':�#���-eS}C����i9��gM> �K����k��<�1�3�(|����L�ǟ��?�Lj�l�~/x��e��D�$k�i�ڗ�S��\z^����%E����RE�E"��Z�ح�Y����]�P�����X얥��g&rW�G(|�.���2xBZ8�<���5�%��$ʊk���&����Q�u���"&ۉ���	������YMbJ��,��G�x+�P+k���S��G�ۯ��8���3�3(}/�bwؤϮl��h
���}�#�{%��M&JzV�li@�!P�$j���*�Sf�K��2���Y��t�L8�2�f8*�>��Y��`�t�`��5����b�cGO���mݩ$(ГهuۺI;�A��^ж@�����0F���Ѷ�!�=E&�T����m���K��xpr��)C@Ԕk0ַ6������*^�}j��z:|?�5{ޝ��-�M}�{R+s�ܶS� �o��/"�{�I])�,}��;�����ȻӼ b~=CR��m���a��zZ)�q��)6\�>k#�G/ܮ���]�aHƧo��ⓚk8n�H�s�������k�����y��4T�qr"� �r��9��6t�x��F�t��Dv���5Ȱ10b�q9�G�Ώ��&jZC]����6������iK��/6�ŋ�Ȯy9���H��-�]��.^��ԓ�A�;��H��Ē��yiD䔖��\��U�1f�C���:��,Ҽ�|�w�)"�?�����2D��P��tC�Q�&;ȿ�ͩdZd�M��f����1����`��n�]�i�	9C���D�בYm���6�(8�
��E�֓�B�n�dB�D����}v?L�	7̶x����L�>Q�>(���ļ4;ͷ���D�g���^زBx�]�7U\����X]A����%�&��~�Q���ԇ&�|˧�B��5���G�y�h�ؿkXNh�1�'�S���n��՝�����G
n4p����4E��l�]��gG5��ۮ*�PD�����6w��*��h���f��=+'gF�Cm�ͪx���+�P�/FZ�9  ����[g��Z�a?��OibpV,�_?�r ��*]�S��>�]2�|9���Dͧv1��g�����:]�m��� ��#�|F�L�n��:��b"�'Xp��~��n�q�(Z`+���K,wU�+���K!�4zL�Y�\����(��,�pp�;��PCV#|y��qd߼��4�	��7b�֍Y��=-�+�R��r��h#R����$~Q�)8})c��]���4�::8�Z���1%Y����qP�㟢u�d!x�J�0����$�ҵ���Z ����[�-=�`O+��s|�^��!w�c ��T�1�ݚ�汊Nb��Ԥ�5QK��h6������DD��}0$���YPkGIc�o���<9�����[����ҟk �f ��D�+�*/K5��.�Dx�-����u[���,,���J�i��kL)�'Rq��3X>�|n߃��*�}���D��h�%�<�*3���e�b��P�=Q}FG�fJ��<�a�NZuF�'Ӑhz�ֻ\ɱs!��Rw�oZ�S���j�H��05d~�����*�߈%�E�6��b~8����w3��0hM�/��^RzC�ť�k���v����2�f�4���@��g�6C%����>��f7����CL0�5{��+[�mOܭXݏ�X�^��;���őz��)�ԼIu,����ȍ���P�ؙ.M� 6�;���V���_��Vic�=�n��FvR���i��Y=�ЊB��+I���$���O�9B�X�<)�������j��_`�u¹�>)+�'����Dֈ9��'��Ab�Xwԣ�֐]����M��HAC��n�����x�GW<�6�)�8�����8��d"�K�v��&r�>��|��:F��B�5�G�#!���~��z�q��.e�[�6�t�����������-<II�u��tM������ԟ�4����hL>Ho<���db�'�T�_�6���IY�=��57�n�x-��ݳ�mQ�v-ؔ���jة�+���-��Kذ�*��������3N�?�4�L� ��s�}T@(���#����)��T�R��|ILe��}�;�O%����� ��sNJ�~��w9����#=ւ��4��^X�pA}k���W{i�P�#k�*fQ��A��@٭]�����z��Bӳ�O�ѡ#09p������+������ՠQ��0��'#_tc��Ec~ܫ�8Ҩ���UHި����h����a��R�<��L-8��*!�)hO��(M}�J�b�Bї0
apƯ����W�ƚ�L���Ԕ8�o>�w¿sm+1�d��q�����|0�
�H���׬�	�����l�"���F���E�O�c��H�p���L@�sl&� @����P������f��5֖�!T�G�R��Z��Ƶ���^-C����T��Z�}U��^l�2��Hq��������z�۝�"&�r4�G"����n��^����f3��Ft�]���v����n۝��MC����9�*O\P�p��q������֭��H�\�-�Qҽ���
�H�n����6�j����B��\�G��
�\fsG:��}\'qc�	�4�z?��J'R�S�M��{3�Aﻣ��c���u1lD#�.e
R�dq�r��<_�[�ן0�9�d��D�2a~�19ی=d$�݄�dp6~��4ˣ�؋}G��"�b�y�SZ��!R�>���ek`� �Ë0O�Ǯ�!(��y�Q,��.��Q�N���q��3�g	2�rM������ 7S�`F̽k��5������ln��R��@��}/�W��;�G�v�qqO��&N�����P˷f�����E:i�GLM~���&=߃��-s�X�i�g��.@��9�� a5� ����L$���Vyy�w�e���S�՞f2~)�F�����(�S����x��9�vO�X���D@U�&�Sg�M����d���+ ��_�Θ�Yv�TY�Z�y���������^��wj{ �?�5���,�C��T|��`�r���{-.���Y�����:yq��N$_-�^(��n�o`ﯯ�Ӣ��6S�!��@��4���E�:�^$�t�J;�f�g�����g���)6j�d ���C� ������s��U�$�O��.--�!~�6l2��8fM*���淭ٮ+pD����v�$o��Z�7�A��7����d� ���O����u�����o�l��ku5��T����G�)*B�˦zM�~x���M̃�X���Y�H�f-�M�\��eq4}��nK�(2MJ��ή�WBC����r�J�P {o���u��j�Fk�l�z�����%�l�
5��.�w�;)u�/F w�ӛ�߂S�+r`�������;Zw4�~�ͳ��?�-~cv�SI��v�!?w��0�����K����z�+Ub���vg����@��ᶣ��/�Ҷ&���p��5;�z>{*ѹ��Rp��v��=���Y�(6FX���^�������%�3��FH$��@�}�!��D��ځ!�Z���0��ծ>tey��P��FόF�ͱ���I^���qQ���Ŏn{�l~�ܟ���s��[��S4�=�[�Kd֍�1u�+����àZa�t>L�h�Z =�𡬰���f���CsǑuF�%�Qb��REr\x�>--@ r�_$�B��Bx�I����5��j�h����j&3�F~�����m
wEI^��h�R�8���9���G�0Ǟ�z��B���I�CT�ك��Wh�p��1$��u�rBlYzX�����%��I��N�M�ҏ-�ޒ?�T�(��ph��+�{b�%�׾�}JY"�ӭ��Qȱɨ�b:�"Jy�`������y9�:��n-������%�P2�'�wiu#����e�?C�_}��b��-C��	�xc�0ߍG�{K"�r����c����fR�v�����d��7z��������o`$-��K-�a�+�{ȡ��Sw� �o*p��<4�vlS�蘶�|��EеP ��8�f�}�0{	��(`k�R�2�s_DSZa��U����D�}e�1��X81|���g_~r���U� ��G��������K?q��e�����Y����at��</�ޑ&X����G���2�5�?�ͦL�R �3�X�i�/���ȟ�kT��m�����iݣ������9�g��9�٫p�
������3�h�	�k�(��������>ksԙI D��NޕNy� �ԣl���Sڣ�iS��oO���^��I:���ť޳�nq���^97y�F�T�-Ǵ�����!�
.��m�7��$pHtW��<I0!Q,(mն���2����c����i��Yx���HEPȬ�J��OOت���'9�z��B��I[0�"�ަ:��F���ƍ`�A�b��R)3S����1�{S@'����-9o����1u���~Tߩ�?�+�۬������7>~2O1�G�m�R�hT
�ufS��e�5�� _o� dd*�nS&���_wM(Yi/\����0 U��r�R���և�ׅCDB�����.@x��B����w�T]��n��(d�ī�I�(��/����g<���S���C���w���l�o�T} ���e*R�Ғ.G�/�5R�o�2 ˸ȏ����]&k�)=���;@�Xb�e��-P������N����2tP�,���r8�(|���<\]�ޅ�e�C��V�?�ރd��M��ZKB�A�N���fp�.M��P�OAX���o�S�.���̏�2��iXtk��4�L�?��]ɤ歃��LK���|�~��b�AM߷��g�'�[�ȡ'��5�e�b4|���Bw�sD�L�б�vX�L>d�4)��O�����/�����yuI��v�b�q��R��'�=�"��\�;�%��j҉�L6k�����ϓ�N�|��DC�u���W�_фW6Sc3b��-BSp�>I��-u�=���3�����!2QB�����j� k	��HF�}:�l����1�\�&/�A��SA��ayҹ��0ᖢ�8O�ƞD�o����b:��	�2*!9'�)OȹKu�y�Z���-z�\�&��y���qȁu�Tg|�EY��W>d2�}�f�ʃ�����$פ�R��>YG��$�)��f�/�����^��/�.�7�~�0&::��7�����P����O�,�u�_����`8W������	���e�I����Ӌ(�}�,�u�y�6[�(jR/؁el⺲n2]`��.n(��[�rX���L1�#���l�QL���8� ��+�5ȣ���fT���@~7�j�RH���w����M��}�,CU�i���Qr#C��Ҹ�0�r�U�Y$�j��hoN��^���:ˍ��0l�lv��x�>�S�����m��>�f���V�t��7T�	a֞�M��U�X���y��r^X2����(vI��ޛ���������$�nA:�[��(��#���k=M��y3�o]�㜽&��`�@ H�	7j�& $#��G���ϥ�Q5T�3�*7<4ø�>�<[��\o����>ћ�N~����vR�����3�0����dD��Ɣ7�9���Y��`�ƈ��z�?���Z�a�y������p��;
yc�Cz�6mg��]ȃ�2�Z�>;�^c���{�o�6d���@^GA�=O����:S�EY�
�uj��*873��y��w��/��E�I:LGԻ�m
��f"dB��K�d.� ��1V�o�C0a�*�`�U�xZa����laNB$�Js$�=0�~bt��kG��͘���hQ6�����*ښպ���S%�����~��La�ՔO[E9�S��gi_$�۩������c�t�5����ԋ�(ږ-T/oA>�F��F�l��Vۊ�O��}�5�w�����^|��̤��W��TEly#���M�ze�(�Zz�|�#�+Fa����q��1v������m�:']&���E�=y>h���@�Y��.~�=�~Kf�͵���"}��֘��n�|Q���-�̈�6��?���[R%��3�'�a���\���4|~��܅zp�X���	<_���{��g�'�A�%�]9�:/5�?��!�k�Z'm�Y�. ,�oY�A�{��p�����a�a�f�S�hL������;1�a����&J����lc0'�`Q��X�j��b�Ʒ�V��H>�'.ϑ지������4���\����e���7U���̞� l ;�YbJ0-�Pp3!�þfJ� ��l���X$B�0�HHq40�}=*5��m�|$���o�;��߫
��KJ��&�q��/!+�\�ֳQ���84^l�i@��W�[�Fo_�z�6Z����$���o��&~���T,<�M�O?����o��zM�R��@WT����cOO"�{1�Q�=��O�۸��J������S���������ݬ:�Vf� �3�M[̷Ƙ��Cb�;��~]ޔ]��yM�3�fE��IT]|�뢨�C��c�����'<��}v�S+~&$� �g�)/����a�����������~�NbT%w��*kg0����7�pb�fx������x/�=� %��i��O�\^Ɉ�w]7ެ*+=a�(q�~Wy����w"O)�:Z��-Bc�s$�Ʌa�����+�+�b�Nq����e��zE�g��p����]+����c� �)QЏ�X��U�\!��_#��Jx����I�`/%����P��{2-�J�:������K>`[Ej4��=���{���_!���{J��kQ�o6�ys�o�¼}�lT�&<I'���^��=���IK�%�X���8�ҍ9��&R]��1��>�'[�&n�殆=W_�ݾ��S���h�넪��j_�	��~���Ѵ$���`	m�$��t��[��B�ۥŭ���ē�́����F'�DvW�bD	A+��� �U�5���*��T�������-�N��+�֥����6��;�H��<TΎ���{|�n+�$�g*��o\�J����?Mu�3!��8p��<�L��	BOM q��bM���.L���M�_/!�Ke�q��,��b ��xӶ� ��E֢�Sc�R�Qn��M4�Ey�_��d\g���h��Z�֚�;9�_��S��� ��C�8��P��F_(_ �/��֝�k=�z�R�Y
���>6q�)#v��nt��Kzyw9�󓓂�d��L��������$�_�ю� r�L�j��$9����t����[���Oԕ��q�"I�'��$��	^]�z�E��3�\����s뾃v� J���v�4���?
�Tv0��q;���͇��d��S�'���'�[lH~��Ɇ��H�zH�5�,�?�U����z��E�����ʐ����kwi�A �; �/��;ϔs%�ȥ�‧X���7�l�DD��j�3��Q:�<������R�r� ���{ި�p;�/P1pF��x�g.s`G�6=G]��<Ą���SP��d�p`~�J�8�)�c,�sj�	�~�!�k����n���(נ�&mz���f��n�N�Y����
@q�N	����T�۹���:'S��A�P?z
X$b	�ȑ��i�8������MU4��5ݨ'�g�dhpN�"��iPP-�Vrܢ'��8,
XΊ)�\,҈W$;�>�ql}�fB��8�l����<1���ڭ��a�p'@�鷣��'��a�(��Y�����y�z������"*�^�t��\˲Daw�B'ʀuaEYԃ<��f��	ȳ�?*�B9 9Cb���\B�RV��rЉ��d�3OD4�����Ɠ�I�$�:\���\h���'�)��?���Z-�7�b��M�ϓ}׌z�V����a���T!֓�P����ڤz�����oJ4R��%����N9�vN��8v�d�����v�U9^�v:�*�Ю�+Ժd�Ra���_�т��zmS� �D{�$����$���Ⅾg���Qj�������5��q ��o�0�������@U�E�#��C����q"=W#��[��Z�A�ژ��$&[dS rF�ͫv|��O*Q"����{.�
ު4�۟��Ɨ7���k?�;`��楣���BE+��GZ��0�^wd'��Y�N� >�.fr1;�����5/ߪu�|�,�e�|��WV�`��<�j(��q�!H����HVq�;
�V�oӱ�Y��>f�^38|���u����Te��]N�2@4r�9�m�]%�C�2^'v�H��X���
C�lev�����şn��є�����c���i���G䨦�"�7���~�6�7+sX��wԍ����\���`����2x��b����*��,�]�1_��s��6�f���f�7�,�$NF6L;�ۀ!S�
و������p~ 7����:v�ǊG������J�3�^!�MΛR��J�2J}���̎�tϝWAʂ�'#?TC�U����&1j`xK�݉	I��.�^�5�'��1�x�ƙٟ�xBj h��LO�&��
�p�O�鲂��tMM^�����d�X����ݧ�$�cN���8iF��}�lo��F�;�`_kM�%є��%u u�-�W�� ��Z��/YCT;3v4�Q2��.L�5S�ɵ����zV���
��ta�{��1�v���qy�N&��Ipke��Ymly�/8F��A�أ� ���h����o�t�K��",dʯC���w����P��)F��e"��R�2���֨�њ����o���g-��h~"z�\��/�w�����D �:��]w.��!��h�4������F�ԃ��I��,.�v<��|��C�[��7ܰ>,��[a��S�����a`XS��;hyb�/�~ 7��> �V����捱�<��぀����հ幝	�%����B1���t�K� �<<�z��oo;��ǅ�:a'k�i��z���$��d�s�Ї�����>��~����Eڡ^�]~��0N�;4q�����l���=������Ny�GSҍ�4^�S�NP�Ҥ6��d��ۭ,kW����;���1��S��"�V  ������\��8���*�c� �O�������~�����
�fz�2�-Q{d�Rm%�������y�������i�t}���	�!fG������c���o�!h�F�|*�`��+\���aܳ��K���:�㸷Clq"�u���`Mv�uo��/f�}�ܺ˓��+I��u�/Y*�(b��ȯ��mf�W�إ{G+ �����F?8���������τL��g�'Qoçݻ(���V���%Zo@�u�|�b��T�;8����j8z���J�bς(+g��G�V3;a?�ʛ���|R-�z-/}��p�8g�֛��*��ۑX��v}��-�7.OG�iJ��E�^�w�����w�䒂��ں������
r�kp�9*פr$hoK�~)fŷ����c)IAk�{m*�����2�1Y�'U�,qi��Ǵ�J�j_͹��~h�<f��3~���߼��-����ʢ�3z\�ڛ팷�|�=�����&�J���e�<�~5�x��%y��Z/Oǂ�ء���ƿ�i/�PJ.�P�uM��kSQ��[#5m�����V��$��'"���ǳ�T��c��ZWv��)U�e�.UW���Xao�Bg^�ba��J�I�����v��@��*��-���7���i
I��ҠDG�=�_��*����k0��R����/ˡ������ͥ�I���lnıI7��(����Z^�W��qϻ�g���XF���|�91��X2l�%�0�"�_��F"��pɎf/����E����X&�D�~�}�����_�RN��C�����h�� ��Hh�Pu�Kƫ�I*�Bu�����|��b����3�v�6�n5�ʛ��]z� ����&�n8�G�I�[:��5ng��(��/Ă�՚BÅrN�~��O��B��}y��d�B�R]��u��կ�|G�p a�$�>o��ᘣ_��q	�*���wk����jO�!�a9�u���\�������5D�E���
b#�u@��1,��� >������k�\9髾��Q�<��/�V�ɘn���%��6>�P�a&��wk�~��;�Z�X{�9q7�����w;a��D'�
�	h|C��*Z���ݼH�aSc/�;���x͝v�.�3������)x�u�So1.�a?��yG�鹪E��,;L����`!/3��n�ҋVd�XOk�?E�F�Jb��K��5��]J`8�����a���Z
L'�T���F]���q)�oj�q��}O��$5kf!�����vC�ю~���iB��c��jV3щ��HŞ������*��\m�P]�O��H=~|�p{
�ۙb\�Ĭ�?�q��b�F�8�� y<)-���m��� ;I���� ��g��{��}�xY�0��t���³�	^�}h,��`�Jd\�Й��d��h����/����>��	�W����bX��k��e�c7�͎����*x�8V2kz#�X��X#Y���掱�ʬg	q�%[��yQ��t�
Gm�s��MC�c6b�MІq�y|7�#�:��Ö$����wp%�~hW v��a���r�E�+�?�D�����(�Є��^�$�樼"�"�M�m�Lgע?�q��dw1!4l�q,��tp�dS��N�c?�������g��~��������Wِ-��M��d0�������]*NQ��9�[Mt')�O27����N�F�6b��/�e�� �3�D���!gH�Q�x^���r���@/��T~����Eq���I!�<IR1z���$4��|�7�Ri�&�X|E��Q?%����[$T���/a1�*B:��e0���;�����w��a�D�І�]Rޞ�3;�Q���K�O���c����R��1@yJn�c���_�tD�qfBno��G~v;�CM��m���h㴿!c�r�Bgo�$����$�WM'urx���bfsެ��;�EςOeE�:�F�Ra�֞a�gA�"RO'��Wo{*��[&m�F�p}�)�_	�y(^W��.� �H�Z�ԯc�)��QI�Ec)Q�,�2��k�TҎ�ym�T#�Aw�q�O����'��k��h�de~����������1W�%`'X~d��{Z2��zץ�Iv�Tdt��w��tc���c;D�'�2���D�����1�8!r�=�
Bհ9����2w�CD=;���+�@��?�&'�Z^�ꍍ 4��-Si!��o��\�'����AH lVh���¦��LŰX�|�M�G�P�*�|�1�p�V�>�R6㉃��4�;#�P�u�p�P�Aco�f��m��n�]��6�2��ۋ��4_�����yg8T
���ho�^I�&���<�C��َ�$�-K˰���ݳڽ��^M�e:����A�-L��*x����E�N�<�ۉ���ՙ./|Cq^�l����7S�BKq-�B�^+���~��>7V�'�Lb���D[�0Ა��P��2�_��ڬ���?lE2��?�g�~���)i�\IqT%�]F�<��3���s�J z`���U�M��J�WD���Sp�e	MFЊ�om��c�G�����y�cϝ텨+��S��s�ݼ��(Y��R�we*�3�Їf��*q���yMOҜ��(] ����@��j�7y��v����]�[�ʇj6�q�)�/Lچ��֒	r���Ře�}C�#&�U���0����U�t�<sP�d�w�"}<�V�������lx7E�e�۩�$�l�g���ֱWD"Z�$��t��%DՓԊz�%�;h%K�M;d}�k��5�ݎ��:��E4XN��~�M�����B���#�g[�Ȼ��'�!ٿ��>+�ѕ~b���@���3'�x��w�q���Z_s����?&�~Ys�>#� �	���T�U�2�䆽���1Aq.[>[hI�q�W��O@�
f�
�(��\��K��QLf�P����0$#0�q�ur[��iZ@�jB%�P����%��e�ڟ'Q��va�Nt�4S��Z(,�q��w�}{L/��������ۆ��Gr��/�{u��'��P�.?V��ŭ�J4EDG\�g�NUU�1(��F{]���$���d�A�m당  FgUx���Uj&'-<��M!~ko~`�M��"%��ʹ��aQ�G����
�]�f�Z�����0f�x�Uq���ր��ں�q�=d�BʆF���r�e�1:F�;Z$s�AS7��?}�Z�\O�{ (�=��qkל��4��o2����ŵLiNgn~��1zr"H���(T��~�S��d!~�g��kC��^b[nd����C��e�k�v��v{��Ө`r�3Т��Vr�;�h��v�Nu�7ׅr����Ho�c�<�} ���.�M�M>�L�᭑=�<غ�){��wЏE��9^�����k�'�r/Z�����A�C��d���"-C�IX�	aG��-��DK�y5�!��.�#���$$[-i�~,�����6o��&%�;c 	����fn$�iy�;�>�5x�k�Ya��	bh���ɦ��&�\k窾�$BQĿҨ�p��B �tho-P���>,v4�z�w�����g�>G�S��r0���uK� ���q���L���t����g6�0���:q Ӡ��k��*�B>"�I|��[GK*�6�
�T�Z��u\��Kf�Twi�7�d��O�F���>ɌŝW�Xbۧvd�����٨�����Z-$n�2
�
-h�3s���{�8	-޽�~�ԙ�D2nz@���iP�eglS����erf�����߷HID釪MR�u�ʙąj�Ue�0���Е�Q8A��ᯧĩ��8j�̏�/�{Q8�&[���(N�� ����J�i�������0�͛�	��?}���Yn�fn��}�x���&�/D�M��.$��|(�e��*6���d3@�E���m&U��(^���y{"�-��'}����fJ��T���U��H*l�kc�gʸtE��u���)��l#I��`M�_��m�!�^����1j,#Sˌyhϕz����r��cq2�SgY����S�+�}�y�P,�Ư�.�r+����k !=`�<k�r�W�-�M�O��[�ڐ�Z:���*�*bV6z	�F��~zo��Bg��N���#�4���0�q-�Lx���G�UV�'>�t�R"�up�&3�r���q�����y��o����f�t�z�	w�;
rs�t��|?ݙ7��*n�i�Q����G*=�0��e��d�=�z����s�Z�7+�|�W%��ۢ+%������I���������� ��)ZD�Ԕ0X �C�	���j6�S4~#�wn���j�������#�BJ,!V� Uܧ�5��|U.�â�-G!�K��W�F�єTC�f���
�͐?����Re��J˓:R���/��=�_��J���v���b�Y���ktaա��q��xd�+#7�tm�K"��1c�����h�����7��@+���o��,���C�R{�|^�lo��=��]_3�Z�����1��������T˞�<x7�(���Ёێ��u�dfWk(q�Tk�Y�	�w�ʴ���
����q�1�1t�\�L�"z�<�{n��6J��'�8�1�n�ǝk�`ŅÔ6>�I7�Wz^���XƯi�WnP�Ns�G��F3�1X`��k�9_�l
V�L2%.�������K���6-B�p��/l���@���c�fJ�Dn|;7N!=���Q��R�Xp$��2fͅ>�� lbg$��33��nx������q�8��Y!���P��aqF;�0�Zlp+V�]
EZ�;C����Cwww��������GO�y�~�3�M�W�V������}��3-���������R��k�@/d�N�DLwE�͈H�sx�����·�l̚�t�L򥋷�4��Q�<��I�g>_w!I����BE[���|ڦ���c Ї��rA�́�����I\����Ϛ�PH��֮]����Ӂ&��`n3�w���E!1H���1� ���#�\ ��`7�S��+E��c��Q�h����.�E�M�����fs�=�-r'B���s3>˼$ȓ�BB!����ܻ��Y�j/o?�Ԉ���ëٷ:	h��+�<���2Yr�5��Y?�n3>���p2A��}z�>K!Pv����&��Z�sH&h�@3��+WV���'�؅�rC�W4ƻ�<�.��j��A)��a�#њ�~�u-R���/�Vt-��9u�\�kk#�?�/m͕�Np�-F v>i�o&�`X�	����c�@�d�yrԱ������Z�����d�-�:�k�w��j^��	��c����'�����f�\�ȿ���h?����{�d��~�k+���G�'��� ��\Hl?wW��r J�#=�K��4�iH"[���~���؝q�fOe��
�����ŗ��b�)um���ڗt[�`{�oڱ�$!��'K����Oa��a�{�d���#������.,�*+��q�1���(�~���(�t�E\�T��S}A,K��ނ�JR���;�PC��;�z�uR�n���]�!�N߮�-��	C������J�c��Y�[k��	�	�����%/}2�Ivde�'o�ߠ����/Y�>�)4޲�~�9�bNt� �K�v�#���<WK�F�z�o��C���z$}��|�R�FͿ����_sq�y���].d�}[�]�נ�@�ƣ�/���pO��F�-Vr~
#�j�/��c����2pSз�����*��5��mI��j�(�j+$���
�'1����U9�?Y��	9�����r�u_�<�~
���� �u<�ѻb�?�pޣ�/@`�qB��s��f:m��q|4�t��EF���?���CL�j���lBn� ��煉��+ټEL��F���ű���2lA��G��$t��j����o`�eSӠ��a�N AW6�ݘ$Q�U�a�S~~�&X@I3���=F��ǩ���]��$���ֶb��������[>����~ֳķ�pxN7=�ꟙ�]�;�j�
7���Q�����P��|�I�gH��Z&��x��u�� �,�1��z��U,��;��(R�à��_�M{J��s��?�/�̣u�,Ϥ���l�7��窌LA��q�S��55�_��3B��y�.( B�DMBk�B�-YC}Q�D�>��e�V6 �uI�0�i����9���Tm0iY�	FO��������t�W|�VW2:����@�F�3�B�ˎ�r|\\��[{�����=l�;J���@�=����zM�v�;�+��-�w< >�����n�fW�(aS�����N��2�C�_�i�� �;�"۵���tz�9�(�PX8�)m��E1��݃1ǆ)��,!��F/D�s-���tE��6���'g���O�$�����X?��=}��/-S��#��E�����o'�:��N�ƣ�k��"�ɟ�6A(_#��_��0�.ӘŁ���39��@oƩ���;��]}x�D�Ӽ\�'����Tp��M��F���n!��uO,���}Q%k�2UQ9�P��%���0��;nRp����ًQYg�5�& �ϣή`�p��,񴲁����'�0�S}��B)ť���t-�� �> *!cqF�k@Z��IU�+ec���X�fї�@���`��]�k��[��Ef
���!��a��ܒ��x����4b�b��N����[\I�~��\�����g>�ցd��� �"k���>9�Q�$X�oK��HM��nD.�3��_@�߳� ���x�ĳq�bo�"!�rjXƌY�GC$��*}��2Fً���\b(/&��F�7 `0F'�A�l���}L>:d7h�Z(@�4S)Q���0r�kz �PM|���a��}�T0�J2~"�Q����95v���t���]�J����i���7�A�|�so��d���|fIg�)�|�0S����.�ۙi��We�si=$	\��.�]B� Psq��4�Up�u	ZO�7�I��5�C{�{��1NK�v�+�m����2OR:�
���:cÝ�K�;A �:a�/�Z6�Eip��Iu�C��r&�+��.�Z�O*��Fܘ�v�o�,l��N�oO�F>�̀Y�v�*�����Zk�&��!^._�����P�����ۜ�3O7 ��w�ڡ�}{s�_�;�������Q��I���Y�IHŬ$X�l"V����RϺ�k%:�?�x+8־[93������H�Ӕ�?
��ۮ��e7���d��gv������d��?��jD�dI���rs��2���� � _��h��i|bn����ߞԽ�J}A�W0?�ۣ0f��i�.��@ӥ4P _��X��r)�)��$�%ej�w�}��%��l�1���R��S}��T;�s��-�i���1Z�Jf�� |�����#Z;JC�Ь[����Ӎ[��`���y��p�<뗻2�����M�<9Q3mW13�,§��*fN�'���T����� [6l��$��o\�әdJ�$���h�L�j"�)����c��J��_��V����C�	�Q6RX�?�<��
^1PS��3��}�˕+<e�w��^G�@��i�Ћؙ��G�����΂P��-�O��dd����_�	���=��qI�CU��㾵0z��ǒ�Qx#��u$䐷`6���&��/�UW�/�mE��:�^��	����F��$W93i0�0{txND����DOL�%		�q�������1�Q���Q�M=4�������#�11�p�y�!A1�T�ݶ��]�b�.��+���ƍ]�J�o�P��bC��l����]-!B$�{�_��~WWpٞ��
�vG4~-�<��C��Gy��.�sk��P�IP�IL�!��U��	:}��3�=�'h��t��6�lj� ��u<KE��4X5��c5�[ǆ#�u_��Fz��c"��,�u�h9֭4�M~#J�f�<�@ғh���iij´K�)ژ@�'���:ͬ�j"���]�ԋ ��*׹��-��f�ȯ	)��q��w�t���_P�:߯�=�?���ܚ��4-��I"�e�%�������u蚤�֟��݃o��N�ͶC�#8��}�J�x����A%.�Bt��Eױ�xy$g���;Ջ�%a���h�`A���$�i¨
���>�=�;��{m>$w���D�^p�,��͚��z��*�/w��w]�\��r�Ӿ�Z\�s1��Kw�x�q~nQ�#�<��uc#'���A=Cj�{?�0p����@1�aʰ�3a[؜���?R[�r��)�w2�8�n̕��D@�j2����BA�6+����f���/WY�����)��T�G�4�$X�叄b��
	�[����J`��H]�~*���` �|^�-����II�)r�h����a�����*&j���p�k���� J�&��í��n�P�Ŋ^�
7�����WʰW����#�4�${�Q�� ��������-s��*�]V�.YO�!}�H 4"�<˵I�/�_�k������O��O�뢥�/:&�QI�1��(���Y'�E_���"SL����3���7��/�b@xF�C���H��!ˋ3-O<�����g��!��+b���)l3o1g�rv�Isqn-� 
����T����:v�F�okɟ��J�ӶS�3�q�@��Du\���:��AN�r��5����L�~#Q�΂r���}3�вc�����Y/�V�Iq���j�؊2YH��o��tUo��=	�3�=��������@'T�����M���I�شB��Db��µ{�$b�<�(̾�?Z��[��\}��X��鞓/�qMQ#YJ7o/ ��Y�n �8��M���ei?t	'�цT�������n1{c,o-n	W��ف�����5�a�Xkc}���"/��;���$lF˓����H����Cͯ'c�Z��7v�$�a�'"\58����{e��9H��jm�ܢ3���p�+2=��RG'�f��-�/��JQO��}*��c�m��嗪So�ۿ�������ly����2�%L>���g.���Y6��x��*�!��_� �̫����y3��)�=|�
L�imR��/�$B�v�Wò�;_����0��޸A�p�w]�]'�}��O(����{?�Ȋ'�y�e4��W��((໣'�GB+t�'�\�e���U��՞��0\���2O6��!���?��-����w���~yr\[ՆUH��~�k^Zf��S���6[]�2QH�@�ҟ�{\жf�i�z�� C�{��[�1�̡m�d�C1�j�y-�u]���Ϊ���ʪ# �G�	������@��Ś���}� ?�J!��<I����6iղ�BB;�~�Ӣ*�B0�U� �L�����o�){,4�ϳj�S�QB���9��F�@Yz[c��	�R����¢�O��!|��7O�^;�����qa�����z��{d)_�x����tg�,'�z�|����QO!�/��e��D���EjX��y*`m`�R�nZ+�ￇ��k�6v'�È}���FW"H�P:p���B�~��&�{Ҡ�4S��߉���6�h�m��I�ı�5�=��,o�m�%����b�Ҹ.��\��ƿq�C4$�T��#���w1{B��.�	�a��hQ-/���9���1�/Xn�L��%m֭mmTU@�|�z�w-|_���� ���'>�ې�1r��ل���mj<Sn���t,})zL��$�G��
RӄT�]r��wq�+�	��.����p���CN���;q��������~�eC�i�|O��L������u��О���������߆1��T�)�;��7ZB�V�.|vh��XG��n \����M�aS���_&D�����"t���IBV<�F��7ֵr��7B���e{}��|0v�7�|�;&ɯIt���6��ѣ���ۏ�b���	�%��������#C��7w�QqX鏯��fa~�ӗS������*��R��=�m^L�vt�;���G���� o��.�_E��ql`��^��ߎ2ԛb�w�2{JY�6��+4ѹ��p0��9�h�o���gx��BE؁��v}�hJ�5��������b'�pt�U�[ �J��lx��A�Q��]5[�"\�!�ϩ<"������q���6v;Tk�5���
+�Ʋ6��-��﹃��:���m�ut��v�u����+���^�$w���_^�#���p_^�Vg�/^$�m��i.6K����"�}��<���ϱH��D�����@g�~�湾���Z�y���@N�J�ˢ���4�n��f�;T�t�E�W���3�g��o��d4w#.O�!���R(���n'(5��B+x)H�� � �i	^}�J;�J�;7�����gUbSk�y�`�8�?��K@�VHE�y�0,|��h���9mP{�7�6��ZT�� !">j<	���a�Qɡm��a�����^�}c�/�ۢ�����%���~5���Wvlo���ǟo�L>l�<=���H�\%����!�!zn2�(�����{�BB�[i&�z޷�c=����ч4*�r��o�Nv��$����Hd�X�V:�T�e����6����i�k��z�g<����@�Վ
ы� ��t�bz��!-��֐���x��������H�W4��>ߎ�'�iϠ$����
�x����ϾL9��l�o|D/s�d�&vF��ItP!<�4�˽���/f���hʛ#��1	���pKeJ��z��R�lv�Ʈ��~���u�[�3eY�lv*���ʟ��U6;�^G�`��bvnE4=l�XB/ҁ���b
������$��[����1`�����˖�`�g�?A<�����q~q��0�wG�x׼Z}?S�\�0W91i^\��Gu��D�ٝ�+yO�MXb�衐M��V���i~�!�;5�a/!�|�c��֪���V����a�&���C���;J:���U�����O!�;��<�0qv;s!�J<�ٖ�t�����1������'��=�P:�q����_��B.����Õ��q�i�yw��]H�,�4��KA��?N�BkzLl2���9D�	w��cx���GK��~P�%
WL5�s�����A8�aDI#��>��?�x��=τ�c�;-����!R��N�S)u6�Oց�y�$��f�wS��g�s��n@׷��a��H^CΰhUW�<��(O�{]�f���~1�����$^�##������y8x�����_�'�HX�� >*ĳ�`�fE#��^��fm&��U���s�	��^.B�`ذWmI;��J�:I��JW������<'�mm����@}�`n�7^3���Z������H�ۉW���kX����;I'EhKq5���c���g>En4�p=�3��U�R�<9���tI�/]O�~�E{烩�(�ػ�x]�n��������T<=�[��z�����(�����[y� X���L�l2��/��H�E��i^,�w�9FHTu���f��)7� � LT��|*ڹ�	�!X�ra�H�� �Xj�Gx�)��.�5YG�a�,�)`��9��wq�b-N����9pc�3(�j����n!F�V�w/� {Sp����i�ߜ���ea��v�W�6Y�~��*�ľ��{�F�2�yY��`ʜ��gC�\��������]4Z̪;��b�"�D�g����}��7���H���h�T���&*�[���S�@u+K+�]�I7b����Vh%�&��=����EƟ��Mw
k,��z��.U�v�2�^7���ĨO'��h���-���e�)�8zX2�t0g�1��疼@P/�h�(�>|�w��:���t��gL��h�R���q�'���V���0���4�t[Amϫ^�D��I��a�HME,���Cg��<�׃�����}0�������7xi�Y1�F4&�68�G�A�3n��P��W�wo���}T�w̄*�@�o�����F�qQ{r
��� P'��e[��m�q�S���� i�هZ_Pg�9SN���?�j�e����WԈ��3fߵ�ki�&�i������8lI,��m��!�S��ߝຬ��;ν+ɩ%��pr2�o\�*$\j~�ǠBΊ0��6^�q��'�2�C���Q�,�%A5uv�3�eyԝT��Ҫ!���{�q�^��������@1[$ؓZH�x�&b�z���.�zi�sg����P���В�����~��oh�e�Y".���gB&�\���N���㠦�Im�����B��Y�Z:�1��s�X�|?��-ݡ�������}L�D���\��#|�����%�Ҿ�I��CQ:�FC�Rm�= +��"ȝge�9qh<���>i�F{�h&V����؈3k!V�����.��uqDh�_��$M���d���9₃;0_��1�E�t�7x�*r'�z������,(�N���(�8�b1�?V���Ɣ���Bv��s �o��C��*K%��X��=�a�Gfdr�ئ��w�LD������h���ͽ�MmH�
��;���h�>�}��1��iF�U���u��3�,+y�yN����>Um�v����k�~��**C�쫞�uk˟��>�+�
#���^{x��֌�?�? �v����З�YV:�N�e<�Q�=�3|����	a(�sofNb�R>�k[�T6+}���39�1ţ���i��pB�[�ëo{@7);�͍/!f.�BI�Ġm=��Q;Ξg �>�ub�;������N�<A��!W��PkS1 ��D�[<6k,i-")KT���`XΆ�[�� o���A�ҹ�5���zy�tJ����#^���b�
B������&?��^;q5��z�0~����AD�u���p|�D��C���,K� ��ɒp�����柏8ܺ�uR�݂֬��"�Ncf��Q�TF �h���,��[�'�v@�YY6��N���G���ZM�^�^GF�6�DZ�';K��Fw��,�K�����7j��Rݬ�dk�=�ݰ�6ȯ���Ή�I��-��9{|��Az��@��}$=�)��).��ziv4���o�x\��4�;N�)TОu;ʝl��$'����3�A[n��k��?�,�uܵ�^?��\��+���W���өҐ������?a����!���$-�LdfiV�����Z	q$�d�s��!M��bX5����}�"W���N\��=O���ʐ��oM�D5�Zg�8�<���pyv�u�q��d�}��:����a��Np(�ԍ�=��ܞY��&D�} ��D�8JO;:���/�p���n�����8&^��%B���A?��|���G|7nLC@u�OR�������� �|`�a�}D��a��|]MOo����EWw��z�������x�����X��;l��7x+��g-���Ζ�ۮMZ�7.L]�u�5ސ�+w�Jr��$�:/���zBʽ��ug���*$���o"aԷ�Ѧ�r�3�N2�6�x�}D����=������\�`�Kex��NF��LG�o�����L�lT(�i��������Vd��w5h�����������[Is
V��A󕩩�����'��*X�O�n�����������⤞�ōxD��[��z�YNXx��\#�G�����	�}�Ybٽ���[�M��̐��c�W���fMt�:	]��q����\�D�iB �-MAa��rR�ܧ�`U9���k>7WKU~f{�q����7�f���J�M�l�/d^,��jQ2�z�<ӛ �� �k��Ç� ���x�췪2�W��ҍ?n����xm!]̺9Y|ms�T�<A��$����?��u�[�U��-�fϊ�Q����]Y�������b����:Q|S
����%�����)^p�?J���O�Z�Y��vfh�*����Y/�:��Yi��Q����<�rrA�RN�tI%'՜9��ѹG���~�&5��+����)�E. �'�$�u#Z��U�'{Uw�?[�±"�9�00�f������H�6��^b�+���Yϭ��T1��d����2�)�Nˎ�o6+vbN�'�|�Cz(�F ط�lz��s|i�̰�8��r�����7��keK�Ѫ��b��+�+sW��-;�UK�n)P���S!�\8ɡܢa�R�X�\8y�8*AȜ����Rf��4/_��"��ۧD�d='?7k��|y�Y�I���<h������qs��������3k�����u�Y�R���<)e���x s86& S���`��}�~r�ˏ��9����V�M)i4���/_e! �Q:+3^������r*��>}�����yy2�2��9�T@y: �h��sS��㶡U��/5g�,.�4�2�m��_�.6��kZ�<�x����ts뿧��RL#஼�/m!�N]
"���w����b�)�_�Ұ573��^���.i�o�^��ܪR�CGU���@���>WOڵޜ5��z:p<����)40�4R[yW�I�d�$-2q��gu7�3=.� ͸�� ��8��-��Ί*��gQ�V�3��0t���q:'���s�Jn�E=Meјpu�$v�����b����k����˘��W.ٶ��hv�u�?e���9E;%k�0J�ѹ�	���z���"�_�$-?��a��dZi@��x_>�=��o\���Wq���ހ��}�~��\<�����m���HM�t��'$KG���⾔>..v,-n�<w�+�I3�||�D=%����'�vŲY��� a&�<�:l�-,$��~�ؚxm�v��"�?�	N!L�/[Tj|w8	nq+Q��ɭ�JK���ķbS��-�}bv��@��Bզ�G�]�ֹ���ڟ��T�[*�"ʾ|p*��)ek�*pX�:��g�w��u�T8+|U��<��W�DU^Z�x�W�T��B�	������=����L*��w��<��{�f�|c�N�_h33>�K��  'A+V��-ˀ��p���_y���9b�/4g�H@����^V�#��F�푲�dG��s@&'�Ҋ��`n#���%�c��yw�哟��2D��dܵ�$S�B�;r�j�|=�Sf��������k�s5p!ǭ�m�딹s���_V����C�����:d'��-������A����8=��mD&TC#�j(�ݒ�-�[K����7�հ�a���0x�_rޫl��b��g����#�ٍ��q���=^v�l ��\��xlff��v]��3�`�����3E6O _S~-U����p�� \�
F�����5�~�c$h[d���#�vn:y��aʴhW�|�*���!4� 	���K��������i�`����;�_�b�����g� F�GT{��+���V����k�V�W�e�<��a�Mt���RU��˛nj���^@Ҟ:b� ���;�POs���b~�/�)�:���.|�9w;hN1�J���$���\z/�rsR�zq�v��>y�j%�7�?<wG��9�p
���L���GJ���л�6�t9!�I�-R/�������_J��}�����Qչ^�Mq�Z>cc��Tz�2X,X�r?���� x�����!�
�ٜ� @�{��,נ;Ѩ0S�`��3R�ǟ <i.�[����>���hV�M��&��8�7����k���
q�6T����K?���h)K�q���$�:-n+, ��M�Bre��S��Y��M���d>�B	�
��ѵ�.�����,P���ǧ%�=OR�g��������->������o��-ll+�䏳��W8��7,f�c^�0�#_L;ef=��mP�l">T�wi#Ɣ�0+�G���؀�QZ�%U.6�z�T�6%@�w<�)>c*���n�}��_�'��,2����������K^uXQ&Y�zO=�_�A`=9�}v��_�xǵ��P>d���㪇+V��)|Ӹ�Ċ'�)OE���ֺRB���4�Ψ�����n<��I��UIBob����3����B��YvW�)�h�真���0#2\H_^&%yl���PH�����齣�t�M>����k�I�}���}=c���e!����i�ĝ���Ȅ�+sa��YKx��o8�O���Ĵg��.�Z�~x��[-p'%e�-��(�5	$���>��%�-Y̺�����r����Ǹ~�/5ʳ�*���-˞Փ����Y��1�Qڝp����/	�� r��7��xX>wz��/<ohl_�=mL4p׺=���{�>;���T]�P�
�"�	��t��~~'<`�x< �3��Jh�,-��y��O�y9@s�h=O�yB k��_�'����ʹw�hʏ�]��f.�4�7�Wn`�WY5�Ih��M|�͕(�+�zF:kud��@��ï"��R�3��\�0<�'Fm����LR�2�����e�tx�~��6.���Nh�tS�*���֫l�J+�����ʊR���I;�`� ��~�XM��ܦ��׹&��1�:���a�|I
&q�u�ʯ���˔��*��2��I�/;*�据4Q�K�oׄ߰9�D�bb�.)�Y�am\��W�]�*1� ��,��#k�nt��PQJrSѕ�,DTB��F�5n�8~\bc4�K���\�|_����.�1�^SՕ
{�V覕7l��B Ip��k�{O\����9������D��A�%I��tp�S��~�c!W�.C�����8
�k}c�������ʄ�GCmc�r��a�W;�T�<*����ɇڑ3��{���4��$@2�G^}�/�o�rC���\����w��������̨������ifH��n��c���!�����c�؁n�+/���d�j�;I����W׭~l�1�Yr8~�xBtY{�03χ�\��Q�m�2���:�؟3��H,�J����Wæ7�rl�3,�1#��w���du��=1w��^���B��;��
�/���|�7�6tЕFL�\�?n�X'�/��ar��Ú�B�_�ᅢ���7+c�����YS������%���ͦ=���VJ�D:�G1�����w쓬6�* ����S��q ]�M�$��&d<�R?��Ǹ}��h>�6B!����Z������s[;H4p�I��������}VF"�λ,l���0t�-���Ď(8�����>�buO/����H���v��iE��KKW�1C.>�X��}�Ґ|g�99 �����-�8���� V�����sl�?��n�Wn��Q��vd`�l�$�<���ۍ�g�R�EU�$T�a}+�ۦ?�U�veH��ΞF$��V=i��$��y�2C]5��)У�f�%��A�,���y��0Z�b�
'�r���0� ��U͸��׶��Ԕ�#�� �WP>�k����1�<{�T
��޽E�����(���8I��#��uD7+���%z����Y(V��[��ę�1 5��l�%ǅ�1ۜ	�cگx��ŕ������]�PFȷ�&o^�e�]F�=��md�K�\	�vÇˎ!њ1��  ���	ή/%�	{�:ө���o[٢Sٴ"}�1A�T���cب�Q��[����]Am�+关h�"_�4$;�=�܅�H��+��}����=a��h��k����ܣ�:�H��<��3�,8�k?6?F��9rו*zA�˔���������7w
r��\Q�]g,YK��'w��߭��<Β���,4������&��)8�B�=>��˷�ܜ"��n��2��I02��~tq�g�{��i6�.C�*��f�x�d��w���F��J��r���VC�r�[[�n�`AKc;�����dw�
�c�1t�jU��'<cQ�mm[�8�G��  g���M;L����|�O��c�Bݣ�����|���Gx�#�?���G�&�������#�"��~ 8+v���붌��̐�+>*���|ܬ��`��׍�w����x�A��j*������n̲+�B�s�?���k�߾6D{��hd�0Y���5Jbz�A+��k4b7��IĊA&�5(~��i�R���2P{��N\ݝ�t�Oh�0	kr��$�	Z�ΒOt�
V���d�Ub,I�������Zʖ����Ax����X�E��ญ�@7}ƀ�x�W!�&�^|���Rp�\�������A�#���e߹���u��I�@_�H.��d�x�asJ�OQ�	�=x�*%~Uo�O�kN@�>J�E� �����,��6����R��ܰ����%�c� ���6�x:��"d�L�h�⤈��W<�J��1�-9cL���⻇m)�&�9�D���t�޲�ac�ဲ���H$��4
$wU�w��;]�����6ڹ��-�%�c�01�6Խ�9bҊ%l���>�4#��S:���� �!�;���-��$@Q��-)�g���DUgF_�C����,ߍ���q�FF��C��[Y�rݨ9½�d�ްn�g�M��ݧ~/;�K�i�m��~�%&_�_|�����1�>��V����o�|Gp��E�`�E�����wgkH\�/�`]mb���Ԥ((G�[n�淞�.B R��,�?�ܟ����'/1�_����(���D$����1�TEꉩ�V�m|�۝��"J���km��~�#EhwM�?�9�N��*a���(|�J]H����U����n�/G� ��O�S�Q*͊_�%�[Ъ��yp�[Z���ؖ?�jd<������_Uޤ�����/���E���R��\P	Vo�;�CK�| M�Re�Q��ϓ�b�Ds�����V#)��w|΍L�s�� ��ܑ҇���+�"��h�_�n+����~��J"O�����j�W�x�Bnc�YE -��]��En���١x0A~�S�{x����& � V�����Q�}�{5A=Iv�o��__�J1z�x�h�Gc.Ða�|yL�7��ɽLbMk4o�]���#O=n|���}�� �W����{���D��  ��s�� �\&�P
�-��v2�ˇS���>��ؿ���:��S��X�F/
e��3�9J������.���J�����4,>0?��g��$�o�5<�������*55Á�&��3<!i���ٷ�3���؇ :�"B3��L5�Y� ����9ۈ95)t.�c��_G�KA�9����R�́jU��;�lG-j[��*m�n�X� d�>:H��rv7P붋���h���,E��͂['��D����$l�t1���+>�L�u��qG���렺mc���
ҿ��� [���|(V"{�i$y"?O��P�-}�oMTW�� ��<�?'	L�#.��t֟�0ju�e�]�2�p���n�I�A&�;%>���Jw�<�N��\����糢7�3����Fܳl��B�΍T��c�w
Lշ��7�Y߀H$6L��1W/#>Mu���O��k^���B�͚�e��Y&�7W�i�-[#�y=�F��%gO��� ~FbY9��nH�U��o���q_p��H��/p�T��Q�\���A�P	H�a����?�&����ԩx�kֿ١�*����?��G:�6�P��~�.@@����E᳠��������8�t.͟2�g���y#��|9ŋ��7��Î�Q�Qޗ���8���d1��=
�J�
/ ��`<ʱ祾��������1k"��ɧ�;"�gWFk�Z�7~��_r����l}�m��.b�0��d��i��3x���'k�	�|}K�1�V�������uG�n	�<4�]AB����*�b@I�̩':ܽ+��KP�C<�~��x�W��_��Ā���?��|T��WY���Et�ʊE�W�ʙ}��r�������<����]�!�|�3����ğ�����
�
۩���b��5��!s��	q
���-�H��@�H<�l����{���2�>}�m�� f<~��|M�7m �8��;�����=���Q�� ������;c�����F�����*5b��,���M�q	!
�OԅgE��Wa�O�;��W�B��T]X��z~M�#t�.�O����返��">&�۟��k)��i	~�6����S[Z2~��DJʚ�_j��Y��Ym�P��T��J�c�}��B�<�~-.n�6n����n�g�?V�<��m��s�)'z��}��uV�Z�_ѧ��4�wr򷟨�:|xG��Q|O��6��y�'s�_��. ��� �
��۞1�~�5n��W���e�hyTI��&A�����8�q���Qֺ�XZs=j:��+����̹h���ː�ڠF+�n�ef��^�=2!~��b���v�g+��JUId����E���0��O~[��l�A��'�;����QM���&�v��^�2͚}���h�������?a���LRV|�L�"�B۹׳�~A;{E�0��g�x}ăy4����n�=��|P��G���4�Z�H�j�E���ã��?Lsm�Ӱ�o�β��!*�k)���LCİ�]s_���ۯNjX/�`qG(���Bv��Z�uOuQ�F��7��+�I/��.b�^[����z�?q�\��e����S�E�7�߸���MZ��s��&����BU�	TC���qጝ/� ���[�x�m��$��k��)%�D�B�=���v{px�N�� ���v�#F��"QaU|����r�q9�1�NHl�r=5�Ζ��=��8ЃV/�[���U�Ǥ�#��6�þ&<S�������^��/n ���_�=6�n�_eыo_��;\�j2pn�)/�T����r���p쐰8���;���Kl�An�/�]wtW?>���J� �Na�9�ɏj�ioQI�C�L��e��͹�s�q�c	^�~�RNY@�����!TT3�4T��� R=������Pb5?�����W��}A��zz��#k��t3�!Q�����x�E=߈��-�G���n�fr`��Ԕ7��(��Dĺ�mp

�oB�7�5@�Y7o7�ã֒����Wģ�\����|��Z��<���ֺԴ,[}X�$-4q�4T�}GW%(��ŁBaW�I����T���G�$����o���.YD$<������S^��_��V�����d!�v^�7F������.�yi1��{���������} lOᇀ�c�7Υ�L	�q\����FϪ�yB-�2��\���"�kቨe1xwM)�	��zYU#�F~���n%lG��N ��:��ˌ���Cd.i'�S1Z��V�c�
=X�dc����W𑻨k���7k�?���v�=*��1��#�-��j����n�J�/�^J�Rܡ��Z�+����wV<h��h�s��|�f20L���Z���N|�6s�$B���z7x��k0"�t�<\E<��yn�O��X��0�ٙ�D�� �0y;�#��U��V�ŹmD�,6����U�k��*���k��9�mH�y!Q7�P5G��Яu��\g��
s�V�դ~M�N���*䀓�7I��Q4�B�"�"ٲu���䚥qG6���:���m��&E��j��1]�if\�}���XD�J��r�@H�o�B�Eұ���U���Qi%5r��e�}h�כg�H�Ω����=X���E�9gH�=F�Ld�v�p�9�T�o��ҽ���5�iwGP�b{�^�5_ XR�;};�a��F��CZB��z|Z�_f��x��6���Rfn-��~�'�)۰��k(p�c�G�5��%�s).��mN�Dq�ٖ��L���~�:�$$���w�#�N�^��ǇM��k7���q<�O<�vB:��p�A�&���Kz���s���>C�����\ӗ��{���*�����o(�.��23�gY��Į(�ѹH}J���s����{��"���ǯbG��M���Rmغ<�BFV1/7��ٍ�bߏ�h����b�T�d�R]8� kA2��v��=�Eh�~���ƴ(+i=v�5;diൕG�D�C��#�y��N��=��;�[?��u�G�����e����{#�G�v�(�ohߢ�>X�,;D2\W�~���3�o��4J��ƒ�(zgb�Wvx%�u��s�@F�*�Le�"���ˈjcQ_�c@�WtXX��=k���lо�Ř>��]S�*{w�Yx�w��Q˧�9� �����b����VeQӴu��zM�(5���̶�y-�ٯ������ov����o��%��7������`8LY_/����뛑̙�.uu�S���WN���a{�6{'N�t]�M�\5�c21_�����A����Y^9sn^��6ӝ4�B�]�nd��"���\��cr�P���c�����%�v�c��-j�5�^��v'�/��i��:�Q�P.�q�zݼX7�Z?o]cy�׈h�B ����Y%���l���a�WK1�N�=`&J��S^�J�9����R�i'͗�1�%�BA�wu T.�{���w�/�ǌ:�c���Wa�Y�5��"[�!������Z(�9���2oF����  I�!�b�ڄ�w�{jҖ�Y�J�k4�;_��g���"�_�[���0}��t���$]䥜�gvx��!���BJB�lNp��b��]��3v`��_��@BWe�3*BFK;��u)�V"4G�`���%-�hu��N�y�3+�~_靨Ο"������,K_п��(kc�}B��K��?�PE%Y�� l���A�V_o���־[�,
�y�TIհ Ēݿ|���/����$�:y"{����Roz�E��� e�BmG�-׿<��w��妹��D��W�*��M�T����'"��Ԛ��/~_��p��������20A�>`l�U�{��͜=�錮o�y��G�U����ߘz�4Ɛ�ʼ��}�ѿ?
3��=�:6���ё�䲧��$�y~��(;�^S��Zs5�+V� ʕ���L�w��+��eG6�Y�5�E���A���� �F���>l嫐�ipL��N���Ӎ塍d��:ְ�ϝ
����ˎ�%rD��H,;U��M�j���j�C��!���j"d�<Ӗ���m� 3��A��z�WC�J2��ߨW�V�<���P隩���g��0����ٶM��n�G�u��sif����S��.����_Q��)_S�#V�4�8ar	��_�z���3�R�躑�fj)��E�Υ��Glr�m�n�ɥ;�rb��q�2s����F�`;:��ش�8�wQ�N��i󮔄LX�%�:��&vx�jS�Y%Z�?p�������� ƚmMVS��jK�e!�4�zW������
 �����P1�)%�3K]�"��,ጱi�ֿ^|����$��V?`��@v$� Q����klD��J����gl��O0x%[�l��m�ш|3�fU{c1�O�qy�)�|�X��=�OH�p?����$���%�b�.���&c��C#ꕙБ��(@��od��;�����,5+�fQ�q$5���[�Du	��Z�2��b��p�;�}�)�bj4?y ��Z�k����&�K�� { �Ë���JQ
c	)�0���9/(��(���̑�:��[��U�c�eyV.9��ꦇ�,[���[�i$����/�x�n)���W5�
I��3�����=��X�c��L%�,PF��C���-���*`�<��eq��R�MW�qv9����df,�8ǽ����ƶ�!�KF��qާ�,�������%I���y}���չ��1��L�$^H!s>"f��w7���%�(c��ٍs~v?0�&UCc�3��b��Ss(�f�>	<�n��>��0�rOV�C����{�O�yB	?���u1����x��{:)~��(ͨ�z~@;ݖhC�~4�`=$ý���ea�捎Ss�Dw�\b,�V��i����J��S�(0��ܖ#Y��uX�tz�j��`g�,�?����H���H
 ���)��-�*8�B-r�*��3��e�E�P5��E�P�j16�[]�p��b`@�>0�\jt�Ӝn</I5yȅi(>�§�ԈG�},�S���� U�#�w>�N����eg1g�lŨ�j�> z.��ԶȰ��k�+��a6K]\Ji����/n��s�����)��5]S�Ε�=���j��
��	���\�2� 3붞L�>\e���tul�Y��1\b�\W4�h��6[���;E:%�����{���Vh'g�=�6Mn9`��)XY�H���Q��E��D/`�M���s��ا�&��X(�rH���Ǿ�C�%�@�Ӹ��H��x�k/R����v,�`e`����~ "��T�1�L��N�����.���B��߯��/q�g0Lξw�kh�<���|"*F_/)	h(��6Di�iȣ��L�#��~(EI�M�Zv)>�g�KZ�]9����p�u��1<//�y1��R��k?5��M^�g(ދ׈
�c/TYj�t֖$�	��v�v�}=�����=��r�O�FYY@E9E*U���?(��&�ڮ{֓v�H�Û��z����]��eaX�($;�^e������{��	|�WЦ~J�L�B墯�{ƯÕ4���q���_��|ҋ�H��H����RG.Lj���"��@�{,�āC���]�S�0@�3�,dh��+�I5�Q������������� �d�蚺��E���ޒ�o�z[���;��Ϧ�&"���_�A������l�m���X�sf���w�T�������۾i<�˴��
�����Zw6t-��\�7E�����L9°����O,aTJ7M�}a��t7����Ŏ��3�NϢ�Z�]�j�:)�׭}~������R6�]֜��Fʝ�{Oy�rw�TI����ļ��ݶ���R���V�y�!�N�MS��=�>6k��ǄYe ���Z�'��5�N�g������y�_����	n���Xo'pJ�vO#�w�Eԋr�ٸN����C5�{������293^�� �oԁ^Y~� @h�7�k1�O�/�w�(�h��ǬQP~����]z�tp��=�-��Ƹ7`��԰n�瀞�����T
͟cu�F�)��*t��` <?��K�<:��r@��c�g�๺�y=	������{wF#�Z�xw�i�t`(�#�O����$dΦ�e�x��i�xm�PpzR���.l+s��g��O+�E�o��{C�hu�v���z�ޑ~"�f�#����U�V�ֲK�n`$uw���-�@�D���r��@-�0��Kl%t��;��N�U��ӆ��;����Io��!2��+��{e���\�`G!j����O� �M*�_��OB����{f���D�2"!e��E��� �7�����R�="fl������{V߂�ɲ�]� yU�S��Y��WhZ0����P^j��7�
��=;.��O0�����jT�;;��/��m+��T�^�o4�	T"�y�6�#j�=!4���4�M>rq-\.�%ӻ�����u�š�����p���J>U_��2�sw])�/0
'�'.�[�U[�1�k�U8�����N[��Clmw��S�	���AJα�ۉ�3�o�\�Pc*�i���-���ɟh'������^�[~ȴ�d��zO�B"|A��S���6�^�g$�M�vp�+ޚ�_,���8�La*T�0�= S�KU��7#�{ԑ7�sIN��`�q��ޜ�?��L�����G¼��wkɯ�Ki�6gF}����/�\7Z�9,�;�3I�������)kتARb&�d���������-�43�x�g�����~>��x�s�8�孰)��ο����lNd:5�V�^~�<�l�����|3Mrl��F��``�#ո�N�u�Vj�2�	�OX#���=ш��lC �`LP5!�W��8 �:RkF��3ч�Y�/��ci-�b��� d:�!���Ֆ��ce����0P������Dԉ�˙
ε��x9S�C<GU?!��u2�s`�Q�?*J�����(Z�5@1�����7d����n k�?�H�Ϣ *+96C���a���!�(�����zd��6��[��B��K���V�9�sG�9h�m��m�{������&�,�B7���k��Y�5��1�V=�Vz��c��_u�-�P���$ �Rg�I���8��#�-��?����B�/�Y�&�!d��J��!u�KR/-�e��oy���A��U+q8ZF�$�tI���D3-��Ԡ������-h���M�o[?������K�r���3��6�#����G�n[�/��bT�W����خ}����SH!������!��9[��|̲U�b�~��4k��W�ҠGD�Y���`C���|��k�7{C�ћ��������Ј�(�:��=��&V�Õ��Ƚ���߃:�4?q����%Kr8�f��4�(e9���Q=o;ʻ6gO�ϑ��Z��Yҵ����dY�<������K�Ak��fZ�g㙢A�ji�Th��kOF��~�).W���w�g;FޣL�H0�?֕�@�J���j�ϑ+����xǸ�MZ�(d��8�(�8��r��N7�+mĒ(��Ww���H$���w&��:l=�~qQ>��\7�<�~!�j+��B�D��%�@\d� a�i-�JSL#������؊ƔEM��"�ES�m\�8�y�N������_�CT~*vZ��g/@wv,UD���N۰b �7��J�󱉦�lR۹���{������X@�9��w�#c�1&�/�3 �X���w�ua�����r)ҵ�������8�1�XB#�gi��]:G����]*d>�����:��d�<��o�N�dU�f���]�Ds���Q������Y\6�h�a��܏x7UT��w�T[+���6�ݒ�������$H�a�ĉ	le!�w���:*l�������`�q֡���&�9ۄ�P�l���?���B�t��I�8xA��Ry)���-�4�|K`e�r��e����_8j,�B��zŀH�y�����2�0ڝ�ާT�E�H�A��`�+7�N�Xi�N&��˔�zL><u�C���JN*u~y��5���3f����.����2�����2Գ�9P�n�
�vU��b8_���(����=�2����0�+�ۧ�%�O��'�=lJ���o�1��H�:_�(��qӺ��t��8�j��,1�z�q�~}�����sd|b��[Y �D��A�o�L����	Hx�p�Ma���k�Cp�^ �b ��A��?�j�e*��i�z��yY�G���4��p1�-��CU��Ly^$=
�������W)�x�$o��,��w�6�,c�H��P������f�~��hD_���)PXE��������P8`��Y�R�0��Ju��������e!a|��߯��Y�%ފ��H��.�Qس�����VcА͜�r䉽�1��2}!�Td*}��.�CV,26Δ��_����"�����9g�q��z��Sa��?`{��8C��P��������QV)k�={�t�� �b�%����V�����a8������=��s�};i�������Qdr�lr����y`�Nc���d&�gd�
�?IOg���ߟ-w�n)r�ٵ��,K�²�MI�B���4rE��e.����;Wn>�A��ȨM�7_R�sk��[���c���X��wm�e������j�.�#Igl�G!��\�^c�WN�x�[�����P�o4�}H	��L�ԁd9�$*������*~����w��ZF��Y��A��I�E�zQ\`V��Hc�E�N��[N؊<|�ON,T���Y�rQ���$����M�9|���U��+�������tIvpkT��'��09��C�&A}bQ�ã��"?��N��������!�}��� h:�:�k��'7 �t�:���u�]�n��N�e�@�+h��W�Q��T��02��%%5��c[�2�Oj�؈z�(Y��Xl�2�Ym�<�-����Ìȸ5��ς��<=n���?G!\񌷿� �C^��rhPJ��.�j�ç��6X0ebE�X�R�ٺ}�A����i����+��{�m�
������r��U,�9ᣠ�Z���o�?]���X)�&+|��B-����6�(��zsc�y�[.���5f�9����Y�^��~�6�D��M��鴶J��mS�y2�ZԢ���=��o�kӬ,q�����a���g͒�qc��3�;Dl}�Ugp泶�L*��H*�R�ER�Lu��H��>��a�%!k���%#-��Q�(�u���a����G�JdDw{�դ2�M/Ǧ��*����G{`���;�5������oӭ�y��\�33���JС�dM?�+Udҁ3c�[5a��
z�8����:mK��Kȿ��@�������l�(�Q����"&RO����Ϯrg(��J�B��4�R��P]�̈���	�m�|��@w��5#���t�fqљ��IߡU��gjRٺ�F����5�5ǥ����9������;����J�_m�6Ow.�Ķ�mijS+�O%;0�����m��Ƹo�·[�Q�+����uL{�Vd�)[j�eA�ɹA�kc�\�v�g��
�2���N=AT�E�A�|zS���8xz����P)���������3(z(��c�)n�ºs��8\.W`������h��7�'x디���b�t���M(/��p.U�}-m��ZT�|��5���.TЬ ��(Ioysጅϋs���Gh:?~H�=��9����x�3��!n�3�o�����Ex�ضc�P�-��@�F�������(���C�fї��Ϡ�< 3�xa��7�u�0Of�8-�xP�ۀ�f����kHۦ.����cM��Ђ0�����������;c�D��*�i��6��9�ka��+)�g��;^#U��J}C$�r�nJ�����x9E�1ݵ�ƥ��d��9&DXgK[h�Z׭�T��03/��X����~��zYb8M�8!N��کHE�F��Sϋ�I(�U����y�a&#h��pUcBY9K���j ݙNm\Q�����?����l����;���E�� �pi��h�z�A��/��f����qpL~�\��x�y�n�LM%���'�\�~т��7�A4嚇�F�v�� |ՠ�k���̌�wHm�um%�""Uj���ӓ>�T��5Y��;MM
G���yq�G�����*b�{�|ګ�|�<#�
͟K=�fiOHb^�;~�Q�G��he�z-�^i��{�N����om�����2,A'�����k�����k�"�
5<�ź��lG��JV� �/����M�1�<����1������xڷ��0I��~�>#|�a���O�TMm��M�{�i-� �hׇ�*�,9l��C)�>��q3xy�@������J[��Y��>�������K�q)��
�?e�ky.s�QQ�6�Vo�iQ�OE5l���nt;ܴ��N�r��I������ƣa��`���ڻw�J8&�I坈��7���{�\F�"�Yʉ0C{�v�.�ׂ_�5�*�* L"�L���鴍E@�}Q�e������!�UL���H��G��2Y�L ��ż=Y���!�w�Ʌ������7l%3]�����\Y����_�K�y�A�PpK��%֐���79��AL_�|���gQ���KJ�F�
�uW\���k�=�R(�GGn��Z,�W4�s�n��6���A�g�a��	#f���i�]�� |�>p{{�W`pl@��XL��vE?п��d6eP�%1N��	�Y��G\��j졓��̱mL�Y�ZO��y���s=׃�+M����p�^o-�Kw#��l�䄳�_9��[ʸ�5J��!��/��Q��%4�r�B��/k����7�B��I�lߚ�ҷ��'լ��t���6����*&ݽ���.���@09�k�d��"8/mdy�p7���U���I!�rO�f�5�"��jX�"<�i���3���#��į>#,�H��AY,�n�����4f8��J�ع4C�{����~�z�� �TԬnVtw��Q�<�m�Q�K^�~ N��lz��疺���>�Y��������8d�k�	��?f��77Jҍ5A�a������C��G��9d3P��?�7�N˿��[j0�BiЬ��$/�f	��M�H�
)=>ن�>�g�r�ѽ4��!	m�$����~��~���X�Khr|��(Ks�
L����_~�HrV*��0��I�`����(>J;B>��7o�El]~^V4�q��Q��4���uЏ�΍]g�6�U�x�Wk+p|ܺ�t��7]@�5�`^rԈ���{�mj�������=Ϥ=������bs����H�
6t&���EUU�Ġ-�E1�} �s��8�G�P�H݋�l�h�^稬H���W'�´	Oy�ձo��!��%��z��<x͝~��JL!����5X*BxaI�X���&_�o�������G��%�6Kt��q�g�f�շ#��K�`�}g:0}�'�A��Ys��b�o���Z$�#�A���ֱ�*����L���ѫR�)�㹑�1��ދ�+�u-��_��liQ�1=�ɳ�C���MD/�A��Ԝ@d��K���Q1��r��4����'��f��������7��Ʊ���ݭ�A&�����e�<�NB@'f�i{PWZX�~��� m;e�>���u���9.	�%�3���!�9�%�d�I��*`�fj��v<6~�vFT:�&|wrTpb%���JY��m���$63dU�����$q��k��#��q(�S,�k��}qbCݾ����t����5��b�}XՑ�BY]�,T,r�O�J��Q�~Hx%��KҶ2��UryTx��#Z\8�8:X�bd���>*��%n�x����E��gk��S�����RDX\W�g�R�(�NG��n-��y�t�&�G,A\!f�5��'�T�3b��<Ӽt��CE���{����kb��4+�ٍg��s�)�{Խ�2��	��������,) V �Ԁ�8
��䏃2<�1
Ι!���Ȇ�'�ۅ*��T*Z��|��b�KJ���M�#]sdq�91�#�:��v=��T��S���ǭ�]R����7�F
�����ȹ�ø�X���v5�F����<�������ˡ��?�]We���2�Z��c��WЍJү2��x��t�o�KĐG�,3g��;k =��C���
$��x�rY�A�L��}OG�.Z���;��.K�A�H�	=��uu���EPL9.p�d���-�}�št'h��fuMn��V:��CV�C��p��$�i��>QY�dj�G�s)<_���Svn���7��k�W3(ԙ$u�y�L�aa��at��m���L/";(���|�kxD��Q-%`�~I��������x�L�����Jǳ�U�����[�SZ�������@�%�F�m�б���\��v<��Z����hSZ遞��.j� ]��]R͸� Y�X`J�`����F�}ĳ�=�_i�v���[=F��.~M\���ϲ���}�ӗ���U_����g��1��U'��3�	e�J��j"�(��fӱE� �n"�ज़�!��r���@]����)>��㏰���~���`۩�Pv��%�X�i���$�@�� �<����[�!k���O.��%��ڑ~
utl+����Y��P�si�-�`һe�dz���U&�ǿ���C}��~�5�-�ѱ}p���_��^y�ё��5�}5��9yC��	�G��� �~ɘH]��t��]���T�U�8I�7v�4#Ҿf<x&`|�}E��Û(�뚇ѦPb!�hJ�1�'^���v�2�ڤ��w��25�8�/��V� �n>�����Τ�A�����X�I�1b�Ն�D<�����f"Q�s����Oq5�P��, �{�{p:¸(�aOM�r �ǈkN`)
���xV�������0<�[�ٙ��\����WlBQ��"��d����Xb4�r�2�����ƕ�ڞ����[�,��#޹{ѵ{q�WC��y�b��?�tȤm`�#�2��'n�m�b?L�K��U��},���R_�J�bu�~'��@�������ⳇ���|�G�#��%S폣�����w�6���Bt�U���H5p���*�߼)�<��U⥯c(�7�!.0<P�M��r�*�JB;yW���o��-F�VM��gh5훴|�ɀ(+�����U�i3bx��K�A�17s�(i���d���b�KO��r�-^�#��b����3��� U�Ҭ��z<?1�  ����ơ�-��Aɳ0�����e�ө�4h��sq�����q�jҊ�O����B�iG�B+���C��/?~[�[|�bi��k=Ra���(o �Z��_����ZR�+*p��I��!�}������y^�jRH=X\�:�3	����
P�v�G��	�˒� ����ls�(ˇ���4��j����:�n���	6��U�UJҸ��H	9�3��>��|M�s�a��IZ�����WͰ,�+;�,D�����x�-כs`�� ={��+.޵�GO�П�:��<z9��S�,��d������|�\ 9BUQ��ħ�6��m�Ӝ�}0;�4��L�ŃF7NM���� -�
 ���W)^�Z*�w�� .�g^Wo9D�F8_�{bl?�:�R��-Tu�f
.�&PH�Kg}��:"M�!�{�2���2�Eh��3��6d([���q�4�vɥ �=����=�٥��.�?�ʆE��e���O��b�|ۜ�lSD�:�,e�K��Gè�_[oC=���J�J���>2$��׉X��;1e�$��#�5�$����mǡ�FL=�["c�Q��:���^d�`���8������tVA�c�=��e8[s.N�̣�y���b��� e
j
L�X|�E�O����;]���u�B{�K'�<�.���<!�{#�͑��:��SS�!��C=?�_+�6�d^�6����z<��z��ɿ�޿�Σ,� �+�ӕP��%���@�~�N��Y!!���[ڬ5/?�mĹ�v_f2������݁�Lﰝ���I��&�5������Brz!>�#n$ic>e��k�|��%��R�T2/������
ß����W��~P�� ��UU{�
�.z)�JG�*5ݾ����X}(��J���P�����D��"1��l(-�G�q����E��~px� ޙ���<F��>HC��z��L Žc���rBH��|qrώ+.�IE���������w��s���:�O[�U�N5Fͧ�Ugفϻ�۩��!��)����3��㴇���t�1�kz�����09*zf<j]��t�82&��yh��Ů-M��1E�yy����s��\Zw�u��?��ۼ� �u�0�(��` s�d�56]�d�����P\m��w��\Ɨ�J�ƴA��Wg7��j*��-����I�{n���p���G)F&��@�D�.����P�~f#SK��:c�HeJn�7��y��ty�y	�\���J��Ш��sQ ������ �	^�yn���wc�0%w2մ�j��Usa[�@KJJp� e�w��ib����f9912x��yA���k4��|K��D��nZV���I�=���Yjn�"O\�?5�@x���DI���kM�5���YͼI�B�ՖF�h&��H�*�6�F�ZqY�޾Ui�>�R����.�-�Iz��.~S[�x��+�yr-�������!��u|x&M�g��a�~ܴC�
��%��l��#J�02i��/� /�ٿ��o���ѷ���.��^�ds��ǔTN�+O�L��F�����ei��mˑ�D������|�u&(D�.��u�{c)<���Bq`4�Л�޷�(%ǁ���N�z>[)L4�/,��rg��Rv�>R! ���n��`��L~�<�U���Fm���:�DJZ5y֔+�t����c��-yև�ԸTv�f�4Y����ik���P�؋ek�7�<��U��%��آ5�,.���|䊼���z��D��v���A�?4M�M#�X�w ~�����y�q7(������l3 �nW���5b׸���\P�?�L�]����լ������w�h����4N��`,�T�ᒯ�L(�ۗ�P�V�X�p�8���|�u&�K��0�g��X&`c��}#�Yd�ժ�zá���+2 �+��h�L\X8[i+�֛���`q�o�D�8���67�_���0���p�=>>�)��C�&g6,�x���������(5�����=���zSR 4hl&F��|���Z:���xlV�#U����!�1�J��.MdJ�oꅳP�K ��q�TI�.ك���+����}frV��
����p��O��#���_%>��Rv+Rx��LG�g/@~�nK��I������Ax�
�&���1�������W��`����G�I4	ʤ@v����hGyz '�MJ��)ґJv(��H7Âc#������c77�sXSy���4S��Y� i�{Q���]���9>�x��� 5�6��ŠC���rS�<��o)�k��S������ѥ[��x̿���e�۹D�%u��C]9ݫ�����P��9�:����=X��G��)���hŢwr<gH	��}h��Ӝa�����7��Mϡ����s�׀��׀<l�!��ЗF�#��d�>jѠ���$}ŕ��j�I�يڝ�j+�"���Y�m�08�k�ݎ�r�?�ro�}m2�5�6�q`�5����?�������L�T�M��J@%MDv̸�+MT�~��3:�ؖ5�J���;K�a�\|_! cW܌+�ގ�W^P����f�p�;.���	^]�����^�
g`��0�}��{]���_^x9�{����~�`�o�UÞI?P%�>���	����(G���#���X� �Md�"����	�����E k��V��Ez-���ܫܯ��<Ǆ�o�gwm��e���N�V��g\+�'��^�8AH �^|@=M<IO;��Wl�Bg�M_�F}3!N�w[E�y=trͱ�h��(<�`B2�����������MS�V��;�Đ������+a-�p������
W��ůL����2��=��C�)�ROT�U�%Nz�r���nEM�l�<�M3���KЉ?ʍ\��P���4�k��s.�"bԵAH�av�?Y�!p�q��@������0
����Xfmb5Pvg��?yHƼ����ܽ�=KF?z�$o�5�Ӕχr~�1y�JrO�<%O+�d�=f0�8;���2҂6��Q�~�����j�xվ�E�h��nfA;���P�w���R����A��z&�S���Ä�~�[FT%�KO|}8��۽���n	�ޤ�޵���������G�
m���NT�mmǣqa����������(���CB?C���Kfq���_݋r���sx�mR�$�Gk��59�0��t��-��S�������y�x����,c��x\%���}�M;�%z���u�����f�1��j��B��݂�9�Æ9���8��7�V;/��c�N]�U4�h��41)�"jn�?�F �is<<�Ap3~,6��������a;�<�ND�y0���i�����ǝ��k�E<�s���p�d�\^�<t�Q��Ծq��kԕC#C)����m��я�L�F��n�����O���v3������=�ݨ��v�8�1}��υ.f�����W�NY� ?��йƏsޜ�i�r�F���� _�� �cA.�=�d�qå�M�+�9��$���I%g$²O������3�יp��o�P��O��?s2�I�n<;�-��7C�^��P�Ớl�!܇�֦� �r����>�b�Y���^	6����؎nn����W�<�<�˱���	N�/��)��\��L^'�&^BA���lAGÝ��CE������Yr�A�-�L,Q���FR��703��Gۍ�!�OG�dB����Ե�>y8�:���g��T�dC�L���c<���b9s2I��5oyٌ1�� ���)[�T�_��bɺGbw�A�pu�8L�O�4XU/��&�!#Y�X��sZ���G;=�%�����K��Ŝp��r��E���#H����2�5����-Ƕ���$<�sat��V�n�?a��J�k�-�g} ^���i�+6B��>�b��/�`'���_˧{���{�h��=��^ذ��/)�=VQq.������>�s��W�Rޭ��5�AQ��a�d����_h>.#y)�#"���t�咯9\0�|!���/5'�!�pa�����5Dgbp��$��ɿ��*�gK{ 0�B����nw��-��"ޢ?�b%�Ah2T�����$n���H�Ǌ�3m���n�����ޥ���w�Dd֣��\}���O���*t'� ?E�"�z�A����ߡM�I��K������gl�'��� �.X�A��r\?����%��Abi�~G֟А%�jK�|G,���%����N/���0QG�9ڣ4�t`b���z'�|K��Jm29�(��.�l�I��ӒZ�#��t�uǭZa�vr�y��۠���Thk�0�� e��Bӆk&��$,gj��d4r�߬�h�Qz����\��-�88gB���n1v�b���B�����8��ٯ?	K��鵠�4��V�'�@Ŧ������=)ҁ���M��\��4.�"�XRl���C`*���Sڅ�1��F��{�U��1FH��I)m��]t�)��c�'=Te���[���&]*�\��2$������&Ǽ�Q��[�Nr@\QbWT}��C�s��I�N�J�!��Yx��������<Y�,z�b^�d���Boߨ�?g�/�O�j=���
�P�S��F��7�MSy3	.���6�I������6��B���U��փ�e�髅>�E�� `���7�`���Il���a���?o@�G�L)���~5dF�q۞Ek3�E$���Z�����F�wS���xxL��Aè<���B�F�x_a0��v����p�yjP��8w �$�۶좴�tW,����Nl�d�l������p�}[��=��m#���a�!W�Ĳ�چ��uN��� ��}�'��e�|:��=Ћ�����;v+9c�g�V�BCS��/�U�`�/��Y{���F��P��Bڂ-��R+��l�^,m�[��&����Ta(pJ�~��2�������
�B���$��{��~hBjCc�Kw�q��$ъ�n��Ze#D�S�[��펦�Z�^k��z#N C�C����&���˔��#j�Xkm�d)|m�y�>
ݽ��P�P�]�0^l�q���]1�?$!%h��8$�#�N�O{J��ף��!��*�;�zM{Ea{��q`�Y3�ɱ�jUU߿�2y^&n��~�� �ȁ�e��h���#��@l�l�Ih_���jmXe��Kp���1���޴��5&�_�Ցw9J��b&R�A�r(�בh�vǻ� t����'O�6���5�z��mxq�%SȂ����H�5��z6�4GZ-;�o�������=<��2	[i���0�)����<�������#�A�u>m�^��u{r*�͚��x�<t?�|4��k ���N�/o��H����L��rY=�~(����G�=wTz����8{�3�e���]�s���5�<��d���f ���dj�O1'�H��#�ڕr�	6]o���Q�95ׂ\���G\4���]3�*������ϳ����gy����!L=����Mh�!�4�4Q�j��s�Ai�>{zR.���T��P�Y^䂦�o���?Wl%{u!
£k�H3Z�*�r�ar1���Yp�g�S`�H<g��$_E�Nt�a�<H/�H1��#Xl�8���\�uT[��?#��58�R��)�wkqww�H)RB���;��C�`��_����g=g�������̼df�$�-���������+q��da��=&�cq��]ꭳ�J�f$�!��>�0t�i�an��צ�eǹ����M���a�mw�{H�KQ�Ɩ�9�" B�g���u���y�[��Z}�N�ͧ�F|*�O3�ܶG1 �W��1]>�xƕ����WV$P��*��-}bJa��q��Y�ap��жy�&��G�Y���}1�z^w��'�Jt�����|����"�f�D�l�W���؀:��Q�WÓ�NW�
�֧ۀ!��G�x�;��UD_)?&�21�+���h]zD?.,G�Z�=�}����p/���P��mOK���b b�q2�_�����7�m�7h���9v?jݭ�0b�@�1@��݊�\��݉|�d�1�aF,27��T�֠��c�'W!mcY�A�fK�-���n{}ޅc��t�*{x��Go�铽��q*~����)�
���o>�p ��=}�oO|�"<�ڤ�nE���;�z�k��"��l�����u;������ ?�����1W��Ѝ,���Z��.�P�q�-B���D[���X��Zс�EW�yMB:��+�'�2�A�_�^�������>04��7�[Sا�D}wN����li��ȾV*��ֆ*1���������k�D$q�� ��AW�י�Ư��E�=��������L*ū�G5��#.��*ڹ��v D囎UC�����" ���ain���5x����8�"�{���N˭��4q_�L��̃�0'A���d)�����������Sv��˩��E�缾>�FG}�=�c5���߽�>y�ڐ�������
�o�]giC_��vO��/��
�|���0�ޮ��߾~�$�����p��e���Rqj��y��SHKPwe�r4�S�0o�ɿ'(��<�0Uuaww���=z�o^�����w2P�Ū�q|ܬ�գ�`����k_��nߠ�X�'�A:g���*Y�1�D��G�/_�g�#sMiV�����!츀�C�W�9Oa�����yHV�7}>�更��������Q)U��n�Ύ�b:b�\?�Ǎ��&�K��¹	d�FMh]/ʍ�qF}z$1���(��č���V�۵��-&u�R+b�l�C���X�Ya�uf�Q�c~��G�&�i�YV���p�� 00+5U6sH�[�&�Q�.���=F�_���!���ރG5)t1�/��G�t�н�������P5�y��<P$�V}B����f#��;�+�d]f'e�,f��a:=�L�����wSxJ�H0_���-�0�zi<l��n�7,��>�\�ͳ�C��e۳��,d{�>�B�h�X������+�9�3�v�w,��Ƈ�d����]_�S�Xz�m��*����n�^���*��_&d]��|�>�Sn�/TЉ��`#�o�����p����{�����qdz���!��b|���E�<��+BM�#U�L8QCC+qyu	���g���+7EQO�Dg��l��A�g����!��A���*L��t�P5dnaE�HY�x|U�����>'��Oh 	�r�n���+��7��G���@�:m^QPF�v�J�3nA��%RC��փ���h�)��ҽ�l���j��Ѽ��(�M4�_�Jڔ7`h?��T�m��z�@!�Zbն1x�F���l"���^k4�l=��	|``9=�b�����������M�dȏЋf����"�ơ��W8��f;�E����߁>�vĳ�=
��l��'O�ހZ{�������m�!���>&&�����aG��ה.iih,�jB3��KJ�W�5I��ip��$n6Cc�s,;w�bwZ���Ă$�(z�3,=��s�ܷ�+��5�~[�:h��\0��9m��ݪ5������?��7&i^8���g��ʎMˡ\�u[�@&��y���N	C2KX�Kj�TS����o�'X�O|��΀����4<D��!����)A��L���S����Kz� ��{�N�K���A�<6�?S��iJ��o���YZ� ��>���c�����>V��&�v����\���ɜ!���\;����C�,cr��������FL�ਜ਼sO(c�Z$�Ez����S�ז������k2��}�y~���^(6��˿�<�R��_��;H�8��4.5�)V������i���1�p�K���O|�^����_/��MFx��^���h�SnR��qY���/,5�*Ƭ��vwԓMV�Ah���޼BLF�� M5�J���L�oW��g�X7������ل�� �yYO�1��B.�썕guHn�s��έ�u��^Ȏ�_�g�7��6����T.�QN`��~��V,��1;��>__c�����W���CW�r"0<�<0�-���\n����D-P����)����U�����QFEz��R�1�$�GJFQW�(�M���E�6�ע[�1�G��j���-��&��ʳ���z,;]��v�y8�f.�cX�w�λ�;K����2�5�y{���5Y������7�/[?����gjT/��&�Ķo�}�E����a����r hRF���c���7��/+�q�����
P��GoZ�t?Z�W�{+��X/��W,�eX-5=���,n�����|3�U�d-K2���K����٭�V����������5Ѻ����Y.�~goOJ��.5��[�JL�R4��{�ҡuQ��]$��%�3lRL�OM,Zsy�ʓ,�9�-���y�_�$PE�Ф���M�,�E�C�7��F����H�I�&��"'�7�߶�������J�H0�%/~�Ý#Sf�n���o���?��7�{i�^��'���wxR��&�}��a�ap�!��B�zYYV��-�Ƣ�݋��<�3���N��0��N�Ӿ���0��kƝ5��b?��F�)ն��g@]��g^���bM��p.JJ'ǅ���1����/����K5��v�q?�k���ꨐڶ���?>Os�|���9��I�Snh��Q;s�}X��%{~`��p(�y�ɇ�g�K�d�X��zӹ~/��ԟ�����|#�͑��U�k[�B>��D�f#� :r��!��r��%��|K�]k&�p�+N�R v���o� ���YAzPQ�l ������_�g¬c��RN4a�c�>f.~�<&z�x���K/肚�3ݥ����8;;�^V��<F��,�4ιcG���c��/�V�	7Rz�:��2��W�ӂ����=.ї��EF������z!X��u'��j�'��3ž��B� 0�i�� �;�9�Ю+9�U����[�g���i;�I�Ε�Ra[�$��_���p~wx�I�2!��PS�Vq��@��B�f_�JwW�)��WfX!��4=��T�8���_���N��OjX_��W,��0Ѥ�g�~�����11�����d�$3���Q��N�Pe&gZt��٤�F:]Ϙ4��) �|��m��Xo��b�xS��&oy����~�{����D���AS���x8|$�7�L�܆�R��2ێ��@d)�Ca��/	�<����Sm��N#��s�W�2!�{޿������z���<�F���q�����f]�="�fERA��O�[,����F]��V�zo�r�٠/�3�a���マ|��s޳|N��8����i��-��������v̎�J�k��O�������c}��Dvc�/Hav���ܹ��oY���\ͤ�=�������ә�}�y���9�F�Ak6r�'9��$�!��˛�2/8��$�z��)�G��6n���M�um �'Vg�����^�P����Є&����oܭ� jX��蜦�c�n!f�S��B��dpX�ܶ-��ǟ�5�������,:ED޳*�?�Y��x��j�i7,"#3���#�%���a5���l����AW�4�mTL�V�%*X�7G�����F�~��_ �ܷS��"�����X�:-hXH�%���.u���d:g}��Mpf�Lʶ��~����h�������〥�e_��J?p�m�&M(�S��F����� R��yi7j4�b�T�;��I�(֎ɱzC���S�� 
�@)�lȎ����{H�1j7���ݯ��}��������4��R��b Xł&�F�l�u��{�"�����x���|}��1���pi�p��)�"�<���ˉ�Hc	kǳ5�QON9��]i���K�G�����E%�J���6��;��nr,� ̊V���q)`?Mh�rxR\�В�7���l�kU���90����#@�~��eD6�yH
6
ss��U�W����Q�f�i��"UW�71T�?��b���5�s�T�FP���q7,V����vpͺ�E�'g9�FF@O7R���M�����ͱ��o��D��QE\5̽ܵ6Dd44�Yv:����Sȗ�o`����0�?&�	,�/e�老f'�)�Z��Co�Ak:k)�D�wOJf�S\)�+�:��~�'ګ�Yql]{Q�;d�d�hc�w�#�4�ωt�<�!�#8*�H���:�Ȩ�G���*���WY[�X��v����jA��Hɹ]���].��n�_d7���i�;�X��3�;����o����Y��mTO������Ro�����|P�XB�K�l���]�d=ӎ� ��/��!��_��Y��!~�-���c���:)��\����Xl�����y'�X`��'����o�=ǆ�ҩQ�m n>f��s"h�}FG�>@s@��Z�ED�W��%��%��~,4n�|�4󳑞E�tWY�_eB������#�Ri�Gg&:�`���� >+u�te}&����[ql�X?�t�m-���9���~)G��n=K���@�F��6\�|G9���_�7���=>�JΏ�w�G�ѱ0`	J���8<?�� �������+�iUr���,�3c��
/�sW�n+�ܗx��ߞ܎�%�e�
XI�d��{݀�A�ϣ�j��� l?�I^��f!����,�d���|��d�e�G�<�VFaC�:~pT�L�L?��-��6�Eh~�2����a�o������J��?'�D�����Xy��Ih<�����B0	��<ڕ��h�"�,L�@��P���/+��s����Ud���N/�u��M�ض+Ke8K��uŰ���)?"�$��,���>����6��ḅYj
�K�6(-��\�6���|��[L	SQ��+2|������Y,ٯf$�A��?����y.����(�N�wdpB�zɐ���ZY���+u��9����Ѩ�����.=�!gy	�}��MP��&���'��g[_�n%�ұlp<)�f���`���n���.�>;-�P R�g�db,=�)f�aq��n�#����<8��gt��rZ�����zV\צ�����c*���B�>5���_���bF �S�1⍇=���������Ck��0}u=`�y�"��s��zldk��XU�����(�~	��@/�ry)ߛC�[ds�s��"��ވ��%�������EKmnB��]��7��R,E+$n+|fB100����Z��5x���³���tP]@]��*u���>Y�X9JR�B���i���p�����&O"��g�$qw�1AcL�_�ܓ�ZƖ��ǯ�hi��Y�Oou ��օ�>�ۤ�j1�nTDi3���'?ͻ���>Q����;�aϋ�+�118�L�MySQ�B���kF�d)�V���֛E&_�<.��_��W0����$G�Q�i�=�8�t�C�X�0�cV�'ap<X�Y�;�,�B�������:�������E�0;Q{FwX]����"p6`���=�1�%޳��ֳI2=.w�����곖%ơ��vFx��{��J�����:��c�G�[(�)L[�I�7A��-�/J�32��|����K�|�c�hL1��^]	m��C�5�u�!�3Iyq�n3�LF%#�8"1Y��z�]V�/����hр���ݛ�sscY��ɝ���4
��V�#�J�����C���x�o��p'�p�jU^�����P��%�H�٣j�/Pg�G�O�m6D�U�5JCkzpv�0>���� i#\fc6���=�n��~��f1��������b��6�efp�m�O�縠Q���&�&Tň��v+��bZ�+�n�	���k���	���_���p���{��}M��A{N�
k�?k��.�D�F�]J,S[���2a�^��+��֘��h����+O���os�{�6og�I�l� lVI�hu#
Շ���_|}>������}��7��;�Jo�'�P��9��x����dO�ІY@q�JX�^d�f���# �.�QNG���p��b�՞SkGv-�ӑ�Ekg8��VN��f������0���������R��1�G֕�u2�6��z��˜Ht~�h^צ���~Yp�zN7sN�;5�hh���Z|�.!����� �L�S�x��l�ܼ��A1D�y�y#d�	r�y6���%���X�tlqO5�J�a�~��e�vz���.(cZЧvP���̚�l��m���� �Ֆ\ �0��(Q\8_���oeaIY�D,ʋ�D��sܪcr*Ҫ��}�%��Nl@{���.�5C<�!��hʴp��@�V�GA�[�*���(��c�?u=�*�)i�!�S��8N����,� ҭ�G��4�B��bj)��F��3Rr�T,q����E�F��䦳?{��u¾x�����k��tS/Ǝn�D7��c�Sit\����tϧTK>�����b&٨�i	�N�[�k1
��SdBC>��.-����9��8Ñ�O��p�8TQC������ 5�T{UVYz�:�J��q|��MmR�|�#8�ыExns���27G ��qX	�]{����� �l��~YÍX�E?��ک�sx�9�=��/q�Zp[��+t�;KF�`�Rz���}+�	)�4��F(	�TrQ7��v�ݓ�'m+8����y4T�CH���8���氄��vq:�2��,$q�J
��7I󂏆6����.�ь�?��5�Z��=��]q2��݄���	�O'f�~������.'�'��I`�&�a)+�^�\��|Y�±���Y�aǶ⬥3��?H:�IV�r�U$v��Ĝp��M����ɶ���B�r� �q���,�;,�H� b����;�>b>�fJ{E��5O���&� �	Dְ��厊��s^S���&YPr��Z�j��'}5�"ċ�0c�{����t�*iZ 44���vl���bwvL�`�	���H���l��<����ck����.����ę����a"j���(�2<����:	���Lᯁ��!A��/�����&��zO*;#(��Ҿ����So.I�|��g�cp侹J�>/��*s�N-G/Y���~)���ϻ}� �>l�N�8��i;��l���Zt���Y0�{Lfh	G�`C�����"2��e�WiIKW��cHsH�ҾNHJ�*�D�:���H2�"A��
����4�#�H}9� F$�����)���5u�^�R��X�R��2���hN�?�(Bu�����ǵm�Q�|c�e,�[	i|�����ٱ��&\z�F3Ae7zL�oe<
S� �}R��?�1�}�:�
 ��MG���\_�s��D�#�KL�okx��ajĮ����e�2A�w� A�t����d�F�6ʪ�Q	����3�z�O���w��d뎉v�������P4T�y����W����-o��0'In��s�s�pE�H���C�����k)t���*����#�{��DQ����t�I�?��d��vw^Pi��O��~�ҡ����T�o[�KW2:<��A��:G��1�i[�ߟ�������a؋��AV��0�F�K͋��8�ǡޞ\�`c)?q�L&�`Yy��i�ws%�\�#1CD��s�զ?��Ӛ�}1��<�pX��UIt���v�g���y+%�S������:a��6��-A+�}\� ��:���%�H�0)�?���f��`�����]�50+9hCY�m����edh32�4�������	�I���v��E���C8g&�S�f�c�ջ���.��v�`�`ջ�,���\��ñ!Kհ��byu�AڭDN��!��d����*�NOk8�a�}^S�{#n��w{:3;�}�ti�a:�X�7G���ߥ����l�&k��g��+�[�į���΋J�E�.X.���w(����Vej�(�v��tf��y�,ZQ���K��R�ד�;�A1#�g��Y���X�9�Pb�d�Ŀ���%`���EͦBnӂ����WE��8����(����8@A����q��ݞ��zqj/!��]�zS�Z:�&`��\��8zp�vV�@�����f��wc�Rv+0ϼ�?4�}]���gzr�^���8��R\��h�����?��g&�fThQ�7�.�>	.�\da�c�8L}�"�YQd\�~d'�ۤG(s��?�t��A����Wn���O��݁}���fп��\��T�y	�K\�3W��L��K}����9�C���p.���܁*����?yP�}G�����C��M���/֫-
z��������k�0w�N/�H���0*�k�O�����%�oJ�S�<24s�œ�&t�)x�C�O���L2���gQÔlv�Ԝ���[�dj��x��:�n�Cctl�Cq���+�����}E�'�q7����:��;������S��K�J�)�Ч/�GH=��d}L� !�%�I��w&(�!D��Iqݔ�nI���"+n����������c�Zf݉(w��V5=#"���?>��,��	��<2yu����G?oj��n�R�E�p'�	�1(ɑ5��Q��'{ߤ6�T�S����		z��5�*yz`}>��z��jVv�f���a���肑�Ԋ[���_*�N;�(�J�r��?Ъ��ސ�:e��np	#�����Em�룸_�8��� qï�L�����w��v/���ē�2�ډ>�����j����\�.1���J,��?`y��ֲId<�{�	S�Ìl�5U|��`,���F1�����A�j���Y�P9 ����v�U�!VJ�i7�-Ir���8�f�B�O5['M�[��ĺ ��@U���X?�m��&&ZN�B8��F ����+_���e^Q���Ʒ;� >NJ6m7���8rP'�RLVuY�V��#z�=wG��^�����C���8O�ZxNUu��}ZԇI�0T+��ܹb��/6�h�4R����4�#f*�Ո��%hC̱R��s�.�kj�_�b���x|�@RM���)�����$����fP�K�ĚS��s=Z?�[���J���'-��[q��q�1?��i�j�|��t��6F	���ic����돫�<��N�B�r��/�&י����^G��<�R_(a�&RǷ��خ7{ȣ���{�}��}.?s�ƅ���vR�H}��L�$5�t�*�����!_yӽk�����f#hTv�Bl�,,�:�n�3�bU�GE/ǅ�]X\���ӗ�2��#��o���ݗi8$�l����b�z�A��8���,X��0�����b�k��z�<u�I��]�?�+O��k�FHjѹ��9~��o`�\�V�x��A7�;A'�VcjRw��Ku#���i�3�*tEY�'���o���7��
1=Ǭ�$��Ɯ5��M10d�܏Ż�|g�Ot��j����������c(|w���s �h��L_ %��b��Xݸ�7��g�f�;�^�~�t�?��u�n����ʘ1��=W5y�xl�>�/��0�+�y��U���gAa+<�
��al��ؕЉ���� ��:P��+�ħzs��{��_��������v��}k�[�A�3��2�((Ց���6�����Yn�sB:2������wzo��
��%yVw��\���$O�/��.w<��O.�]��I^��mL�&�}�m�`ڳ�QE�<.8z�M���OH*�ߊ�&�Y��D���=�Qd����O��d�:�>�W��
{�ZF��{Ē� 
V#�w�
Dߴ�	���D��Y��UT�
����0)"BN���V�聑�^|����d��O�B��k��U�WpH�<Aӆʝ����2�V
\r0r�/�udʐmT�tG��T�[k
��F�%ªnc�m=��3ǹ���*��Ց�vEl�{�#K��B�n��J�K�UVR�����F����sW�1���/X vzT������a�it�-r�Hy���R�tS	?N��d�'��ټR�g��m�z>Ũ��~��ӀlB�\��S�a ��fp��|h�)>LJ3['³����k;���X6'߈��)�q~o���
����/���
�k&�-�n6�[��y��,�VW���ҮF6��g��B�A@E�⏗hք�En1���f������ Pww��e�f=���jsݍ�췇JL���J���=΍e����ю��X�	Wy�q|�.�����]�{񪮺ݶ�
�
S8./�0�Zw�g6���x��&v����m�1���Y_�6��j">n��p*W�H SA"���^M(H�=>�[��:�"h�1�!�Y�>}믤lA\���W�Bn�L�H�nhlWSL<���<-�޻_��}���y�����!�[�?蔐�c�i���qa2h�~��ϯ_� �g}�+O��J�b�Cզ�K��'633Nd|s`���&�
��$S�E����V�Ƶ�U��t�(���n��4y6􌘳���[�nt���r�p�2A̖	�-��so<�Q�e�g��w5�����2������Ck�%��*D<�[�:��Z��v��=����F,u{���N�f,  �� ��9g�ءG��<ß��^���yo�G���� Ɓ�
��P�mw�MO�eN�CaKǠ�9���p;��	�0�H2s�������ܺ-*�A���>��߄�R )REz��bX�T��׆��2"5���*��N��EA�Q��$;��t�<�T��d�x�M�n��f��)�s�Nd���6���/k��c��j��I1����z�W���!ŏF����.�Z{ԇ�����!�v��9ie������}:��..NL�:;T69�t|�ۼjgeh�xaB�ӄ�Ζ>U��;�s���'@��;�����Ve���ꇘ�rN����#�HF9�kB�̬֡<h5�A��D@R����/���Q�l�`�⁢�4n��bt�#3�%t�&h��B��s�2y�ܐBL��U��U��[���2�陿;��
��b#�PYsL�[�^�iË�����P��v4@:��9	?9��T��9(,���f�AN�oPB�j~��z+a������o��9��M���Ge�̛�|��<D�h��"K�����I�A��� �gKH�4�ړ�N���/e��0�F��4��m��47��Z�"�@ ��.M���@���{NlVN�r���9��Z�O�W\<3ȢCe/e��B�}K�?8�ƌ�[�
��o-O)m~8ǁxc$8���67+���U���v�YLr�R���Y��J��s��ab�����r�@�&�)"}4�)�Y
�#U��tg��d���h���5�g?�_Yܧ�#�l�i�h��3X��0�6��'�mR9�z��;�XH�s<ks.0XNf,t�	�H�흃���R{��R���g���:�������w~�_c�^��bI{'u���g�~?8~�Jv��6��)ԡP�����)�W��X*I3���i�oA�5�/�����x�6cýI{_Lg������.ş��y���Gw[~E����#2x�yn���s�D[�/>�%�k�i="�E����E�m\�����%i;�r�Z#� �،�X�S�J~&ǳ7{Fp�Z:1�k1Y�d��-`ݿ�nV��� �!��ʼ61Z!z�9�(|����Ī���O*�H-$��HIɓ�������4���8"Wg�i��j-5�k�����c�<H��P^���z[6w��x9��\�5�m�sJ��"�R��m�yS����N�kJ �FI)+w}��������=Ep��FP��Foe'|�l��.嬳X~T��c[����e����XܣV���IUN��؝�H81F�e�؛�g�a+����k�[ǫ+���h���CCs��%���p��_%�Ѩ�����Ĕ�щ4.h�s'��a�,�����Ceq`���k���nC)��D�&B�n'o������pa{c�nw�����M��5
��͔�07��c��*d'�����ϳ̢��<���a�@՝\�C���Í2G+BQ4V�ߎ�?�?WQ�a�O��*�^�;�P\j:��q�T�	~��s��
�[D��k�~��գ��'թ��̮%�9�[Nd�j\Ȏ	X"QuW�l��5��9��yk+��Va�}�D�\����*�J) ?��oOG����lhջ��m�0l]?��
R��XEG$����x�gޗ2�k���<1ӧ筪F|J���δ8�Jb�.$������ѳ��2l�?2�\�k��6�����`�	��qEG����9�X%�7����V
�-qu29TМ��˃�;��>n�RMI3q����'�]�q�(����i�� g-��%,@v��) ��- ����cUs� ^�gj�#�3�nw����[<IR�b��w�֊�m�@���T��g-���3�忖cEW����Jh��z4R,s�\䴐�������6m��V�/u����6�R���_�0D=���U�y�;*E�xz�9Az�j�k�_Vk�P��l]C
J&�1Z
�V5���>�<��Ǆ�����UmM�ӏ5j�	����$���D�:>�=S]������B	|��8�G�1��v\�ߒ�/f���m\x�տ�M��¦w9T���~��8'F�b^Y��W�(h�Gqbg{���@����2�f79�K*H�w�}����w��,�������~Q_�UJA<���3�d]-)��fs���t���i	Z�*�E_s�K�^��`�z��&�F,ܫ��X�#>����#�-��,Q�b��3�io���|!�[��JDD�j���@�	p�ߋnP�9zo�B&��ƗV������{ϿۊE%(��è�Hl,��Y������>�_��Y��8��c᳂�ѝjm��pݥfb�����ԡ����WF�Զy=S��E�M�5�D���h�|Q��ԯ�v?�U���D��RO2!R-�m�%V�~ֶ�����<׍��K���7;Ҟ�LUX�JJ�2q`��ӊ6r�U|j9ӧJ�^e#=t�`a�;7�y�|��m�=�d�5ڔ��JjiXF�>�z?!��G�S�'HG֠�H$-p�+�V_l7:=�Su4r�E�w-s ��Pc��gzn^C�Zw9��=����gE�H����8�:��m@�g�֪�6Ɏ�>֛z��(V_��e�|�N��jvc�[Ǡ�ϼ��W)� ��ؓ�����M?R(�$�>�rT?9��Gh�兩F�QҲ�J0�x�"�l�o��l�w�M��h�	�|��)��/��縥@J�rDyi���؍���T0ך���c�g�[���OƏ�,�t(�k����P� s͖���c��Ղ�9T��Ol����%�;dh��R� ����l���M��4%�7J�w����b�]�� ��UMpx"��r�@��e�g��V�x�,��[f`}�Dp�	��L�"�jX�vV�EQ�$�1����}C
�[�_�G ���/�eѕ/W���_Ds6�7;��V��9�2���{">`�4k�2uj�a�~4�0�v�Ҩ5uYf.S`��B�� �|�]��u��ў�G����@�w8���s�>
HAs�Ʊ�|bhe���A��\���񑈘2�Z������B�7�N��bV
0Q�J��:�;�m0^�����&�[��{q+Z;;�!FMJB�%q-oZJ$������E�Yu��f
��Evm�V�ܣ@�N�z�2��*y�.3e̺��I��m�qV�>���@��Z�]98p]ؑ��a�v�k�h>��'H��̈���;mq����tF'8u�嘎e,���b�_֑�ҩE��i#�Q�o��f�v+Q�[d��8�o <�u�%͈�1��v�,�U���Si Ю�0�"�	X7�Y�Mb�����J\Z�Ap����a��p�R�2�]�ݍ-�!݈�Z��M�������v?���Nr8`>V_'��P&60#HvX��l:������>3u��e�)E�"�^�R�6�8�%?�.>�?�B�j�$~|:�a�*U0�#2�o5�z1jԿ�fQ�����喱:buu�B��0-L��+�U�P�s����R?��==�T�z1Y�u�B���4�p�"�
2VQ�`o4��0����x�gkeeA.��M��S�Qq�Y\�n��1~��W&e����Z*xr�.�(�F��p&8 zFg�����$��9�k�{��J�ZyRA���:@ޚ�����\o��m�\L?y͋�(0|�H�NvX7�?�����듀V<֣��ʷ��(!�ʃI��Abny޽m\��"�����۠E6��Ȉ�����b�*�5WЌl����v �����S����5>����l�?�<T�{GK���������VA�B�L$S�9��z���2����E�Y �bR�4�(����#�
A�er[�ЬW�h&���Wl���< 9t���W�i�3^���W=9�o�Qa�@k��Y[���ZHa��@�i��*V*�KӒ��Fk����da^��ݲ���a���꽘���ا�͵V���TC^�iv�{F�e7#�CkF�ΔG��S�$k3�a�s�W�ū�b����o^`.��m��*N|*Fo���^n!L�A�����S:{���6�0�+�����՝DXCn�W���H4CD��˟&�q�X#�3�L ��ѻL�����]5+���@�K���V$/���Z��9��=�<�	�D0��U%����f��������ą�:.p>�]2�u5�����Ub�#�1r�yE�e��V@��.���?Ct�֋�a�W&�ȏ?>�z{I g��s�
���+�*S�~�2�]i4���s
co&E6�Lr+�ξ~��bن[��m۞�[�q�ʥ���W���Cu��F�gZ>-�% �&�I��g:��lS ���H)���ؽ��^�����p��}Zx���o�����;mu\�����j[����q��H��.j��&�z��SЋ.��U����v,Dk�!�p�WYs�3�G��<Sj�֜5\_h�H3]C,���Q�Um�kћX�1w���?�K�-y7i��Y?�%�"����eLe���K�
�{өe��E�A�8�[(O�&�G��p�d~]����Ia*ӱ���Xm���t8�E��44T��=�t���y���Hq�2��fJG5�(cJvZm���<g��5CU22=���O^�<���8,�3�N%�f���_�n�b�͍�Ҝ�3W*i��-��I�Duc�V�PB����'�C��ځ0�h=��Cf��D�^Y���2({��ć��荕*�A��+�YJ�C������ԨR��m��[� ���� �1�L���y��=��[G���5l�{�v�r��f�x�	�������V,��m-�Q�G��ƍ��!�+zNR��i�#�1Xﻕ�b)8��4d1�UԨ�4nWp���K�rg{!�i��qǱӈhb|�޴qW������L��'P��h���$��+��~�?�cU��:��h)��������86"a���_�@��z���tM�d�8{��&W���h������.1�9*�*�-�	�{)H^/�@&���N~eLM�m����*��&��F�����984�3!�	~�"H�/�*ge��dN(_㬢�t�[G���N�0��C�lD)���X �kS�V���+�ta�\H��Đ���*t4ϟ����_�m9��]�F=�B�o�jL8x)����
7���p��Y !w�@뵐kIS��
Lk���F�/�#]�6�`���{|�t'X��r$�\���g��G�:z�_����&�j|����(ր�朌��ĵ.x%�_5�Xvz�b+00P���?�ozkY��"���nv���"��R��������QC��~�ѩ[$^*I�F������6'֮�_�UZd��vg���>����3!SSfC�
��*��h�����uÑ�#�i�/���3����y�!�����=�����I�H�2��|�Ӝ�68iqd�J!�;UQ��Wq���z�MO�I	Ͼ����|���+;����z�ߝ<n����ܛ}�)�>��Ͻ����ǒI����L���<$�ɩ�gc�c�"ۤ%[R5y�kj�<��/)�H�уG���T���Y���������<�Q�"!��(�0Z<�Y�A�}�֚�����w%�2z�U� �"�cA��FK"uf����KYj��u��swI�6�P�;٣E��I�����i73
9X�7���zl�c?��ԝ��+5c	n���i=ޥ8�S��{�����f��.r��|�q�pb����V������j�k�Gq).��)^ܡ@���+ŭ��;Ŋ(R܃��Hp,8������?�X,��'sf��=3��Ü�tK��f��q�#Y��8^�^ƙ�!�g��	}xޛ�[���P�f烷ֽ�>�Kا�N�����#nOc_����ͣz�����! F�����U��;�ɵ�ͳ�%��)�Yi�<���A����O�q��x��ڎsKM���/NLG{��j�8g����x��~<.���q�I��!��Ǐ��q2��&�{����C�$7�H���.<���:�U�������$SK��H����z�<ml��:�0j)�g�̚&�����dԼݢJ��''�"в�g2s�$�������0uas.�ZNѩBM>�����-sD"��Ik��BLv�N���^j����wX<ƭ��R/����m1�����8X?�p���c���b�i ���>c��l��9����T�__��1z��@�0!x�3�?Yc�%����� ݜ����WO��iD5p�wtc�	H��tA��c�ػ��꘯� ��ף�f�.�h��k��]��?@%,��w�![{�v����jŚ��I+�yl�.k/gD��*�y��r�]a��&�ы�o��
�SZy��.��N��v�1���<��|��5�Ѝ���fszVz�{-5$����WT�2S�%>�MV*���ݯ�"޳QC�@Gx���<��;�tO��x![4z:<Q=@���4�N}z ���y���IZ#�%������(;"��ᮔ����!-��S�T!�I��iY�,8��*�&ꥦ{hY�{Ep/��i�P��hM{���.�S��W_�(
�"���r��V=��wc��w�E3�y�ڠ���{D�X1}Y(Yj;5�����<oҽ*�Zev�Q��c^�5ѱ�����]���,Y���� v�"��1�t�Z�e�~u��Ja'�k��ح���W¯h�q�6Gz�H���C"E�=�`��<�k�5��z#���hr�z�ln��Fp=����8��O �7m����-��EI����@�����~���@f��𸗭�+%�|����fXr�s�S���=(D�rcQw�Z�!S�h�uH��~`����|�߅`�b<������}ȫ��	|��2IyGӉC���~�0�#Q��U��1�P����=Z�)51���J󖞮����8i-�쥃��:��p��5�5S��=x#��h��}�/�:*���l����z<_���f�G ��/$+���_�~�,`��k����`<ǎr����T��~��mG��tš���S0zn��p(���#�w��� ��ɫ��J�Os�ǚ��e���0�&�����i��sz��Vs?��Mw����7X%�5m�D�,�u�2�^�b�ى���EB�LXǺ�:E&�.�-Ƥ�mW5!�sR� 5�M���5�%~��ƕ�����n,FwŠF5������u_��:	�<���S��^�@�<�`��NN����tXR�x�I�t���p�.�1��d_D�K'�`ǥ��/�����9�?MP.w��u��H%���4��,VF]�򦂹��NQ��$�}����{�f�~��I_k��r.��<����*����#�/���<�Cs]�����B���������4wF�g�P��P�l9�Px"*y;�+�d:r5�O��d�gn*}A���o����KB����;��4d|e�.*�|����=}L�vb� M�I��u �sp�����;P^WmϽt�&�KL&d��x��{�ZWk�5ʼ@��+	����qݶ%k�d���:<��F�>c�4������#��R4���֪|1��CMַA�T$l���p�z����5i����U��n�_.fk;s��W�.� ��6br�S��y*#B�9B��z�,�QV�����Ũ�l��/>�����a��?�}�Fy��O�j��Y�&K������˨B�4��zk�9�s��B8a�'?����f|����dZn���H�G];e�F��'�&Udp@�(ͣ�"��LP��v��a�_�~?��`������W�v��b��.�;���$���}�+ΣŵA�-Xĥ&!+��%B���%�68����\1����)�Ë��ɞr���~�%1z<�K���J:꾽�	���9�����q�Yl��cH$�\��%�݃5&8�rg�����H{�]�P�_�O��b����uQ��b��f5��3Xy%��"��"a'l�2�����ܗs�-n-T3#��C���ֆ'����J�Z.�B�ō��oB9�a�h���s�}X�a8v��Us86�"|�2��}n�����)�c�\?�75�|����/:��\J2�����=av��sϫ��_�UV�����̸��䤵����}oQK+&g�bV�պX�18�J:��W�C��`<��W0N:�����*��7�v�q���b��W��e��� =m����x��|;#��M�H��<�M����`�uɎ���*��[E��苤��YΊ�X�8i���T⏧�����-�1��P���ȷ�C���s�_?u���%<5�="�������p�Į��qa�1����G:g��:�s�s̬V��!&�o)��I 7�^�ɵ���c�c$�@E\F��Z ���-E���C�X��g��׭e�3|Ve6#�0%)�|��|�$Xk��鈟3b�)�ex?`p.|�����V�H��������.R�oV=<+���cϧ�=��ү�{���~F�gb�8�*��Q�����z�O˕�`��?/�Ŭ�Nb�o���m��6�p�(0������D�ڹ� �,g�F�Q2���D���T2�uÿ�U_�V�ĵ*O�Ì�8�Aϸ�.�Z��_�R�6���m����?}^�X|�uЇ��4�.�z�-�݈d�8���n�3=	�p��Mo��o-��U�V�!����'W[��a��a�=��P\�ז~z𹷞�z���ձU"�0�ܠ��b9Q[�c ��о_���9h�w�ˬ����h��O��*�����(Z��wj���>yG=>UR���s����?���tp�Q��̭�p� �[����YWR���๞nݿx���ܥ͓h?�3�`�$k#KCo��R�P����3�}Jy���eJy�u��ж��nѿ��.��_X�Z`�Lp�����L����9����r�V�/R�ͨe��QՂ����"�zMY�����F't�X���4�m�O,Z��=�T�	eB������G��`�����j������V��X^�z�9?�׽������{������hw+��s~���8��q����cܻ�aV���c�橨��Z���X��^y��#���R֭�q%w��$]�Sq��ʥUk�GiW��q�i�4N����o`�C�a|�1�Z��N����l�VJ���1^��<2�`�ͅg��)~�2���)��|�9G�,\7A���T+���˾�Nb��:��I�,ꐲW�F����>9Π�w��
��5�h���Ö�ߥ0���i�����7�9�@�B>y���$��K�f.��A�4��R�_<`q{�����w����
�Z�hg�F oD�L� ��}lw���q�Piګ��m� �@���w�j|CWNW.Ff�=?�J�n�L1̜C5�Qҕ�)�L���P�L���>�/!���`߂�/i-�r5���{	�_M-���UWn&tڪ�{N0�{^����A����$�&�|�mǌ&��;��cky��,B�h����������/� ����y�F"�g!ϣ�O�1�����w��\�)ˈL�A��K�z��-��`[*Q��o�~���L��#*�܅L���Hn��h�+��j|\��~J -�*��u�#Kk	CD���W7�o%��2�W${J���Rir��Ϗ�ρQ�V��?�:�}h�&m��E�R׮}��0l�w�k���������j�Ct��P�U3��-^
`\ǧ@�/�J}�-�`C���g�^s��a�=��锈�^L������x��j�m�GM�� 6���veU»��t�)�<�:�~� ދN���=E�?5��|�������g<H���o�}"���lsn?��2M'�,T�Lj�*�KZ(������Qk�_�4o��T���� ͭ��]��4݌��t�������߭����I��sC��d���s�+����D{2��h q�1��|���t��?���1��g ����_T{�+��&�%�>�T䳄����b#���}�¿�E��W�"�ʜ	`R���Y|� �%+\�&In"p5��`��_���E�i�&X�] ��(��l�5p�v2$2����1��B�zq��C�Bʨٽf�pE��l�,�}��z�qR�6��)v����VF�=q��?�k����k��$�S��:�D� �o!��n�{�Q�c���)[<�!�S>�_�h��)��kZ��~�Ńs�3HțȂi���?˼�DR���P�\D��0�Z�nj;���:���	}�>`�̽Đ�g&�|a�����A�[g��FSċ��z��|Z�;�A���җox�һY#ݤ�Q~!ufy�Sg�8��e����{�oV�#.ش��2�4�v��j5�p����U<`2jx�W���EsT��j���/�f����{��ת3��������M��Ċ��<g��� �B=L5C��4��+m8���~��7Gʖ��{��5QO� f.n��X�Nx<��	ѫ�I��� ��%��]'��,��]��J
f.m��5�}{��s~��h��[��V-7�/���G;� �;l�@����I��п�0�[w ��#tgw��&��U�k�s�A��6z�b*ujy����>�YQu}��s�:��ϻ���B���J��`:�α7�g���;g����Z4ϳI��k���,�󫬂�o������V�_�I_�[;n�O�g.&Ǉ-v��qJ�E�g��a�� ���t���ҫ�����h���?��K]�^�⯠z�ԏ"�[#.m�v�H�����$f}ȏ�N8��C�:M%h�31���*w�<o�s�)�����K��@G�2�g�fx?����~��Fo�Q���s�~���2�*��P�O��ُ=P4���x�c�P��0�݄Px��@Op15�>g*��!h#�L�t���`�gz��uڳ�2��/�ޯ�~'���|��$�ZAfd?�w�@�"�«!���^ua�\3C59~��p2�J�!h�I���8q	+�x%��\��������rd+s���A�_��3OĈWׇ�����dmW?��z(羋�#כ �T�H��\��E�&�+�K��Je,��81ĿԜ}5�u����~�i�z�I?`�߻��{�L`��T�6ܴ�Ξ��0�C jq\�B9!��D��/V��l¯&W�1��D�3��;8�tsN{n'�{��^��{�G��}��wr��}/D�����q��%[�J���Oz��fީǰ�eF��^l���)6D6�#!4<��:س��l�y~��~Q�����ON���ӿ9���V�WY�����B����
C�d��g)�P�r>�%���&$�N�zCH	&��BOpGe�sθN罎:�n��0��j3������x�XZ����G�~?���5b>Q��ӽ��;P����*@�n;*�Q��gϴ����8W�<�_ax.ɀ��3�m�a�������Z�v� ��r���&V���S�$�Z���Ӡ!�c�W$�'�t�ⴺ+��Z&����4���׍�Ar��W�J�z�X��L6��^1>�t����4��C���3esW ā��R
G��Ӷ�k3��nRq� ��P*�������WVr5���V�O�7)���yk�+�����sy>��iѿ�7��ĿK�
�6t���Kj5I���c^�F�U���zv+%�/�6���:�94�co�+�>ϊ�3��hZl�cB]IHnv��8-מ9˼�����1��T��eݛ8�y��eX~��>θMw�en�?͍�`�y9b�Xc��"|�`�����1'��1K������D���5H����ĀU1���\՞xj��g��'v=�>�;zȟx�~�>��8���Ƹm%j�j*�twI�~���enV4/(�_|h��Kz>�~����x�
8�8�j@l��=7���Q]�%ɣ~�5�����K>̫��B�֕�d���Սה�3>��9��FČ�Q>��-��o���{'�z���PM�\�˪� ���Q��U�e:�ڀm����^Wϵ��.o�מ�����'|�*e��]X�֟� �j�o��!��ˁC�Z/�J�Fe;9\�#jGy��7���=�#���GY�G�S�����Lԟ%h:/���R|�g��%i�ǩ�Q.w)�������!Q���#�%	��y���CN[���� S�ޝTS)Y��� �K�����b��&P� 3�<�����i}K��qjt�����PD�&G��	�VE��|�[�&� p/��H�J���GG�}�)��pe&o�.�������?n���<���b�K��I�ɛ1�zd\�������&��\���Ӻ��k�F	�	����{���9�c��g�:�-ǐ��#4�^�+q��z��,Q�[\+�л�M�C�M���XXpV4%��?�bTҼ�ఙ�0��Ⴀ��
�!� �J!\u�ٟԋ�K���j�u��Qw��e����2w��^�8{�¯�ƚ��@J3'}~�{g�@ݵu��2{��8-uu�3Ӱ�Ͱ���E�����'§;���F��$%:_d�w��8���sD�A�i���Ht.�Z����a^��2��q�7m��j�N�UΫ�Pc��ԓɥ��4���b��=��C4����'�\��8�C�Z�N���k샴��r�ң!k�����~@^���=�^+*�!�?f�c��f�8�u�[�(���$b;	��E<�U��ư�X��4��A������n�۲Zz�������qC�%d:v���D?B�lH�[1�����Ե�ǽ�6z ����#���O~�={�CԘ��F�b8J�z���}	��;V�lN���<���1�8]�OJ���i_*�xl��K���%�����P���ˀ�'�0����A[F�>�P�thl"_j�^�5��d�@��%kS��N���*3��s�˵�g�U���u�L�Zf&g���������W��ѢM p3p����4��=����W��`�ea	C.��og��<-��nV^�L�KA�
*Y��z��9��y���T</��㗜��R^j�~5HO�ѣc�����S&�}���+As$�QFk�8o�j[[�K�<��ǳz���#��^]߀W�!^�dC�m��"��}��o��=�m!��)��7]��.����b?�Ex���%ͫ]@ս�4OC�k����Q��#Ղaf�l��j�����i���r[f㻱4f��o\R�,C/�<���K�'�6��C,'G��Q5
�z�.D�r�1���H�QoS���bєP-�u�%�o���������iX����]c9gTB��~A�8����l�p�z��s:H����g��#]-��WP�Џ�0�L��u�~��'����!�*�4d��'���\̏�"��(���~��\��tuQ<�8�l@|���<ʖϼ�Ur�i�Z�zC:D�Ѩ��̰``����!>F5
���0zX����X��s����U�,��;bE2�ep�m
m.���BE	�*s��y�?��%R�	�uG;rK�!���7 ܵ���XQ��*5� ������Ab���SY�';k�2l۽��m�/����\��7�`p@*%[�X��
�i�zQ��E�6��Ùe.&$����#�W������"�y�h=�����c	�E7.,�r��0�WU�Du�� 9��x4��Ll/���=_�u�<�P"Z'�7��z�ľ�SdW�uA�J8�|��G���u{�r~L��N�0�ю7$,z0ٷy�G@�[)�,I-�y�%����s�����$��ˆ���	��t줢l�Ƃ�S����LHGn��`�7;�?�jN���X+��:�����0O��B�;9�3�� �-�ubA��Dĕ=0�y�aD��m��q�.��1$(1�����;�aU ��-Fm�Lo^E,�9d����u�4U>3���e,m�i�W����Bȴ9������tH35���s82ѫ�w�IгY0��Ƌ�b׸���y���{�R�!�]hY��?�c���j%x��ɢ�X��qd�~�}2$Y��~�Ve
��I��̙
���1>���?��_���p�h�N�Э�lV1�$P}>��u��j�A����<�P5 g0�yKsb���{��ΥB�0�g�G�Ф�f��d�% )��#�{��+�e��w�:���(�J�M��[�µ@�tY����ĕ��ٵ�ֲcpT���F�{D4@�s�� ��˔>�P���	��.$�@.�P���6*�
��amS]��5Ϲ+���|��� -�:�p�`C�F���Ke��,���w�|
�9��`�r��;��5�j�j�v�:�n���9Ȉ;</`��ޯ���������=�7��;����U���~e�!E�Q�*.�N��H�Cn��@�D��_>���7���N�~/+�t��.�Jg��Op�Y�U��d�$Ҫ�]��{m]�	{/zߚ���~C��]u����-�E�wX�C@NH�#���xPz�H�OW"5tW	:]?4�B�/�#V)��6D�l�������k���A5F|�3O�Y��w$t#����۷�n�&�cz���xk�4�X.�GR�%O�>|�%��qt1��m8Z�����غl2}}Ard��+\P��y�8Rg��仇��9H���� �TB"&�q��?��E�����I�������d�>�r����ۘ�8�7X��:~s�R#���8 �m�B��Ï㸛D�ш%��^�������b&리&[����o]P�锜Q���X���Y���jZ��# ��=��E�/�Hu��3�N�%�e��}q�V������r GY���Z�GV��_� �pS�)I���Ed!�^�r3C����pX���t��G�A�rN �;����Y�"l�`#��KT{�!�� ����YEq��v0y�;��*�_F��7M.��	�{Ӫ��)�B$p���]n�\4>�_o��a��=�6~�ZY�`!���L�0h)��n�4�\8w5����:�mb�z\�ӆv�;�'cIYzt^P9[7�f�zѷ��͢?9d�o���Øqf��v�{\9O	+�{fb���T�����^��R���s��Lp����t֢s�����V���",`���ޏ��Q�'Y4T�5���N{`�,�����=@��~*�{JL������7\>�ye)9�M��%q��0RAI�.o؜�v�l���P+����bbK�X@eh��,0�6��,rr��Tvs���補��jA�:�V����"#qCy�?V7�a	�q\��Ez~�|P6�>Y�e� n��hx!�c8���S�+>i�=)�T����oof��W��W
:����}-��њ̪���w�0F�-�h�Wp�5����?�%I�0�R�?J���FW����	�}��ۡD��gR��dC���d�P=�Z�G�H�����'Ҏ3���H歎��&�5)���D����m�-������uqa��!�:���,���?8��E9O/$�A�hXgMݸ_�� ��{���OŽdퟫ�6]+����_��`�+ŇA�{w��j���⏡��x�sG����;��"�qCّ���(_#��DِG'���Z��*�t�ؚ
Mf�Q�3ڴO<�fw��x�"kBΔE���JQ ��Kk���FB/�L�>��&���#��e�o���uܼg��������,��ݢc(��x��pp���(���R?Kﱟ L���	������5�p��C�Wu��1��Yj+�'��)�ca�l�9�?��zne��C���ֱ��y���@��ue�)�����k��r�y�q~��ReE²� 8B�<����<������ܵ1��p/�\�	HY)=��.~�>��D���k뀈��Ӱ��t�q�٩���-�揼za��G��'�V����5������;����H�h3OVY��/>	�1!5ȅXńo\Z��Ё��KNI�Zƕ(�*.����#��r�� �J�t4��L�2��;����W��5h}�p��%����f���R��ʀd����I�&R���š��V�ɀ�5
e)����(M��W{�Z=�*�	7,�g�o�ĵ��yI��ʝ��i�p��-�B�bܶ&��ɰUw�2��']k�	I"�W�H+�f�v��Q(��E��'У!�%�Y��x�K��y�k�F%�EO>?&P�ٹ>�[�c�a�Jdp�ܓ,�zm������+�3��[h�p?��w�1�}ں��o�d����_Ы�"G?���N��D� #�ȸ
ʈ#D?L�R+�m�Z���o�K;�*9C��"m�ƻm)!E�V���mv:-}�ĘeT,rZFHeq׫Β�n)�b}Ǻ&zD�k>(����̫��x�c����d����370 �i����S�	ě9��!��~/8��x_�����Z���7=LC�r��1��%�<�c 6�*�3]�)��6~[9Uw+��`"�ZĬ�8������ɦ,+�JM�髚t�i˱�dC��m�_���o	��_o���p�h_Î�3�j�g�g�AX+S5�<^/�3�;0�2�(]�\��y��q�<��O�� ����o1,h:|EB���Q����o�] �8��ݐ�U�k���Mm������!����>f4m^��0E���.�����E�P��Iυ�q�Yq�Y{�?�9�lb�L�H~l!�f	c�e^;9L���rR$�K#N� ��'�+E�LT��$O�݅�S�ppH{�gw	��Q#nB4���!\�F6�F6y�Dp�M�`���Og���S�0���E��:�<1���۱Nx����g��(��GmK$��z�&Do�u�w(����%��EĈ^ܒ��J�����^s��G}�ZWU��,1�9�)��'rpG��g�)MH{E��t�Ʊ��j��{���
X�Q�Tx(�����?S�����=�{bt��BkS��?�M:�7���-���k�T��a:���|'��B���G_>���鏔�ob���u���)+��R�D�fꑅ���&��Y �Z8L	L�>b���<�y>�("v�@�W��ќ�Z>�0���@�.R�āc�C�	uW�k�p0d��=,��\�U��I��?�LR��CR�tŃ�υ�m>�zs<�X�`���^�\Kxq]�3�-TEG��L�q�a��y��k� 8�_�w��,���V҅::EIz��]rm��Eπ
�B���ӟ�.K�v{*������=�6�i���q.C_������ߠ#�2���"^csg������3�K'�sE:�vi��bO+��il���,J�n>����M#W�>'�U�y��P}U�y�N�m�B�Q�����2��K�{,s��Vd���ƴlC�w�-�8n>�3DSPN���?��
^Y2�og�xqz�d戲��]�if��f�o�!����N�+�.Nժ���H!�������<�ڟZR^g�A�D�?�[M>}�.��ș�17tF���u����"q9��Մ��k��5�ި�i�]�=�q:<g�\������	�j6���@���U����c�
`z����%�ݷ<�EΠH��~�%n�'���J�{�v�0�v�Wٻ�:"�Qh�e��̼'�]��=�M��������n��-ޏ\E/�V�����Q�I	2d������t}�8au�z"��.��,� (`x�y��5�ϰ�����Z_���r*-K������<����rq���>��|p���������Zj����ƥ����e|<�tG'�maH<��o��ۄh�"'��6�{O�����U�^'څ�W�����Ǻ;_ݻ��B� ��0	��Ow��O� Yl��ǳ�Ɍ��x�9d��l�`�\6
\�{��@���m�XR~�ӑ��{Y���U���ҿX�r��Ϗ���C�]m{������T��&*J+8�|Jn�͌@��ϸ;'����x'k�u'2};(pIᏼdl�M)�YE~1;�%��� [?�"����d�7���w_\��,oK+�m_I)�Ԍ]JFD.V��<�
I��u�E�!��p�?�{����Z׽A�VS?n{������e��43���*!��� 0`�RS��a���𣚻}�]�2A�=����w*\s�U��HfR2�y�K8��X~,�Iҩ�T#Z6��Y�k��S���U{4���Ɍ��ޤR��~J�M��NS�`��.����i����W#���� KsI��s�^}�ռ72����������xU�`�T��b�2c��78����2�bmy��2��2z����=����bs�i�ޱ��f�t~�k��޹�L�ӘJ��)%�|+�����,�ݥ�/a�.�G6
)�C}�޲|G�ز)�R����kf>&Ew:��}�<��O����m-\��y]��������i��z�l���H�/<���4߼�p��&���m=�`]���-�R��0T�~{���"1:���-)
A���3e{�1Gz� ��,2��u~�7f� ��gX����Q�,���{��4p�	��a�R�������-��Mt ���f�ĝ�r�h�[n�!*;�inn4
��R괸K>�
�|��v���R��U�x�?݁�����A�%��&�d&�(ğ��_+r���Z��)�G�@r���H�<T��B�h�{KhY8t�RcLҍj�-�G�HsLp��[
��ѺF�H8�n[��Խ[�٭��=	@�|_�9�����H�8#66
��]h�F8!�H�'R��ƺV��z�OT�UKT��23��W�P���-�����U;f�
=�k�:�M���$m�lAdP"u��u��ۍo���f��*i&5�sٳ,|����ǲ���������)=�ȕfw������'��pw-Z1�Fg	�}�M0�E�Y����0�I~l$1� &�#@8��;���Xy�wq��p�i��ta���Ӻ���V_�ݺ;��ꀤ{��+�ɢ��x�V+�`d!�d�G3Ꮍy�X��'���M��ϋ�ʂ��c��>�;�$j|� �|r���M������$�Z{��"��`G�I�S���Ώc�u�@������2��/i�v��T�w}�G�k<�!��F�����I^�chO^�ϥ���P������{C5+�7�3�e��0��bla��p5�Ϋ��ZR�����<~�`����h-�S:p;դt_p��RUf<1�blB�ďP�5\������*�����F7\�rh���~a�>jey�u#�zJl"�ڠ&����J.ɠ��.�=�Pg��3h�cU�����y��ZQn��[},��[Ӳ��1Ղ[��ZO=���(ahu���*��A���uҀ�k�I���BW�ǉ=���RaQ����!23���B�G���Uf^܌���F���5�	��"���U�������R�N(�=%�������f�EB�/k�^XU�%�L�+~dϏG����@=�3w�3�7�i^eK�k�s�@�$�YDdvѡ��5��g�lL���%���EVG#���O>.�s�i�,����:p(�r���[�}��y`�^ß�#ap�ǳ<�V�ysE���`�b�b��ħȶ���1T��B]��H��*j% ��鯨�(�so;�����'���*�M5 V�(0h(ϓ�P2�/�}�}[�7��B�!�[��+W�����t<����ֺ���nq�a�f��,�u�{�������zl8�Ǔ��eƴ�oȐ�����j�髆��c� >�E���uZX�1R ���C)˫���	�5�&\kQ΋
����������-?J[ P>�7�`�.�\O�"y������z�n16�&��U9���mH��������x7��q������j( Ӹ=�_MJu��,���nG+�)!��֙G��|=�w�-��R00����;�l�s���
X
�-�ǎ����`+T*��푷y��/?FM�A�F��Q�.�+����%�g�G��r6�닚#��{{��X#�Mt�,���k��AEƠб�Cx4}����B���C��s�.L�[6L�2Ӈ��k��6�k�k+(�i_��֟Į�(�G{]V|����`8W����"��+����e�Qp�YՅ��v����}32�Nܵ?�2����Q�>���Z.@�������f�+ׇ���R�6t�:e��EUA��,���I[����N��C�\����B�r�����r&\�2��o{�qz�I�Qi�b#�C��C��+e�u\����%Г�p��IbmI��$�V$���1�`j�i�_���ω����&<.{��(+}�8�잢���]��ڋ���VbwL'd�uv"C~�wrq2Hw���'��t4UJ�z-d��K\�Em�zm��[
�@�%R�xB��|+bq�q�Z����'�����K��Y��]���_��:�;��+��[�6����|�����_�I8�RZZ�O��5>�ӿ��m�ͺ�U�� �:툨�����ɒ-��j�(�'O{��d4-�gY�2��e����?.i��e	޵�(��mבQ��.˼��rH�dB>��>��sB:n
��[�2^��s�GA��*2���/"�6̀@D�N㵥j����r�������m��i��8@,����ǭ���k���fwK�o�?I��P{��KB:T���������ǻ�s:B�~~�Ε���L�}ۼjU�[x��:�
�J�O:��!�N�jm:�}�p���\���Q��CP�-�Y5T&�O��H^�n�88��I�Em�|�9n�AfD���Wi�7�P�w$#�Ѝ�t�I�Jb��u�4o>~�de[v���{a �
aƍ��� �B�sq�}�.�&$.x��@ÓȥgkU����<�@�����"��1Zn�1���9�48Q�@�@�ۉ�����S����;��#�Y{S�?�q��['GF��ɾ������7%��p3Q���͢�-�������!ެH���P��H�ͤ�o�+qz�߮�����6�c6ت���`�N��l��𠶦j�nH�Ns�	��^��e#��(i��BX��mx�E�2��-���T���U���&���E�>��٤�چ]��B��u%O�ˮ�(�:f����a�H������NDVڬ�N�Ͱ����;�Eת;E��O����X�w����-��Wc܊]-�q�%���7n��\r�Vp��\/�U��t}kd
����!�g�.�9������u>m��V��(���ߺ�c� �5w�jҟ���}�o%y�[��}*�SS��N�uG��H���,���,ƺ5����7����/z�js��sv��xQ��*�D2�ѿ~t�n�x��-�	\���Al]� v�4���p�s�D4�j��7}�zy<������^&Xp�e�s<(H�qH<�b���E~�8P��#�S�G�� �y;�#�^��{1L�~�z*x�s��Pz��CJ³�\�y�V����5��8�$���j*��m��cV�� �#�7�B(*򸿳R�D��(q.���K�'y�uZ�:F�!p��Ӡ�2��M6[���70@v�҅�&v;�14x�����I��۩�Yg�����Pw*'�<���~�n-	E]M��1�F!O�X�S����4���wt�����x'r?D��`�C�NEzX�6_�r��R;0�9����^A.�T[QOp| }D)�/w�u}\������.�"<1�% �g'M�=%�q�B�J�ut���E����Z�S4�1�����&��0lj�>�L}�Gw��
]���3�Bsiy��, �4~�	-�遅���U�h������[.DHC}N��\a3K�94ͺ���)$�M�_ݪ����@n�ޛv�c�YKi�+R��e�Eͳ!{'�~m��kf����=(�����s�:�j��*�$D;=��Z�4˰ȿ�V*m{�X�
}�'d}�Y7�~yn{���*q-`�V���
���[�����֢��q\�v�OW�5��Y�j}�?5��Y:O��
��y~��5�T�����L����� iÚ��L�����v�t��;�r��QF�_o��f�1��>�U&Z�0X�bB���ˈd�ʹ7�[�\a��5�� Шg.98.$���K��4���T��3�[,Kt��o��<K//�!�3����0�
!�a|��C���+� f���Qf�;kM�Lj)��ȫ��	��R{/3~�u��0[��� +��\Kî�֙�*._����6�1�=0��;���
�Pw��t$T��+��ؿ
�߮K�����
����mi������[��FZ�n��i�t�n�7��}�9￯�k�����~��1�<��b\�#$��|�Ja���h=vi�[!���N�SwMہc�4���P�F_���yK~P&�e�c%L��Ҵ)�ŋE�e�5Ɓ�_�Ĺ2B�'��f����g�^��G�Ao�d�y���"�oj9�4W��Y��YI����g�(2��:��L����o@�XD@�㗳�J<T�t!�u�Z��p:*/��z)�P�����~��zЍ�%��]���8�C��OD hB'z˧a��Ҿ~ִͺh�5+�3���nb��C�ÿ�\c�BR飼��Q,�_GۺE|��Kc���sv���ǮXk�_0�j��bD����q��q��]��~�F~Uݯ�K-\Ƨz�*�C�5nN}H�Ղ��Ɵ�磔���e
�ͳ$hi�2S���9^���gw�q	~�.�E��	n�v��'�z��$�.�a��ϓ�LL`��k�^Q����������H(�^ٔ�м�W�������E~�ɽ!�(:�"�����`�~��D��	�Ġ���{%�;b$+܉���µԦ8%�.IL�j�O�H���(J.ۯ%����?Me?�������h�u!�����s՞o8�9H�-dT5utЉ嗞D;��(���Jy6u�b����J8Lӑ����I�￯�r�쏺�IC��N3���׏�|�xc�Q��`�
�n�6�H��Eid�`|���*��	[6��)d�`����� ���+��{���F��|�><�B����6W���~�%y�ȱRn�n +����^?a�p�`� �f��q�&�D��ݥ3;�9?B�*z�Q��}m�k��H�������C�51!��=��v�g�xcj�{Xhy7�< �Zfg��ڗIk�\e�e���\Z�������=e^9r!#q�7d%��鷊��!k��
K��B���63�°��r{��r��+��g�������$y�ʱ[�^8�."�s��_�`!�ЇI�����,��Uô�=��dH�r��e�����M�3km^�h%gB�yAB7�ɰ��-�2tt:�U��ݬ�io��}u�+�����Nh��o073Q�R�I	P��ḃq�z�$��d���В��q�Ey`=�RHs/q�S՛W�K�dAƈ�K�uM�T��"��kJ8��� �:��9��_�>�K{�u"�fA���]S%�%|�Q٥���s���������u�ml�rݱ��Qo"Jy|�1BR��[�F�<�ݭ��cΚ��d<M���P�?~�
�����������u?uH3�RR�ѯH҂ϱ�Y�H{�JMI!Y#�����<sD�n�N���!Ѳs�� ��~{��ԖP��a~��q>k�������ts�� �^L�ZJ���'���Ĭ�;�[xIk�yP���"�U|�L_��o�Q�=b�Lm�D^�Er{���U,u۷BR���'�_�W��3�+$���
�b:����zirf���)��-�$�!:O��Z���yc��k��C�1g������W�Ԍ�����
7�
Igng��G���=~��O�#m�j��~f��o�8l#���B~}���� PE�~���J���c�tӴ_Od����
��VU���q���O���C�ܨ`�{��*H�E����:�^��淪 Ey����˩�4�Wh��s.
rx�4+x}�΢yq�E<r���;�9�Ec���{�
:	�e���ᚺ<|;(q�Ӽ������O%�[��gbbI ^�Rnn�"�H+�o�Ƌ�� �h�N�~�yN4vh
+	�[�l�jn�q�wP8֗��s�E:��A</�����lcZT=�F�g�/�<�KL��͟�1׸���W�qt���o��s�I����Icg��RY}ʝ5�ɉ�/�d\m�౉�~#��b��=��s�;��G��bwE��FZϝ�*��o�����Tq���~=Ͻ�Dd�/l�k�k1�u�c����<no���1�y��]��,��N�~PzJ<��$�A7k����S�W�c-�]9�B�:��=�K<!�^���*��C������ۋwZ/iˇ�갘e#J��3�(��Ny, ��u��NH��L�K��}��Ў��s'/�GS'�*�O�p��K��A/�S3(�Xé�5����M��4";��eƽ��E�8VD.Mɏʶ4k����2?}Ɐ���Ĵ��LR�M�*��z�f�b2��Jp��VI'2����q�gP2�������@`!��	W�k/{�4�0���,z�.��s�W�e�f7Y���ƭ��T�p�Z�i��^p�r-+�L���cC�8Bc��d����	�ͷ�	�.t��Tbp���C�{Ӹ�g��16���n���[ -\'����)O�� k�h�/��������Q"���?�9~�����+G�9�8�9��@��^`񤸆@9M��~G����-�x2ߝ��ը�����X�ё#���Y�ƾ|{�#������ҍ��LH�O
�'�aW7Ե嗆���،5�~s��<t�i���0���C���ֺ
:�y�,?�<�k��+��Lh�#s��,��o�m6%�2e�
rǵsmҩ?t���j]�Ax��e��;�s��Ʉ�$26y�1S�u�q>1ML���w`�n(l"T� ���<�W�7(������r�$^0l+ �`kD��JL��@63������]�{� �[���
}ު)T�6W7�=�J�E�D`OQ}u�K��7�������J6>�Zxd`IԋI�=ӊ\� ?����~���1�'��aϐE��r���O#\�ܰ�F_���|�F`z����|,Vx�u=I��[M�W%��ա��#�����-��Y���C��\$�$S��x;ڬ����o���u��Q���Ap	fI �~�5�����A:���n����o�7_��o;��3�Y�=����+� ��1�����U:�4�H����'+�N����C�Y܈R��:j�Gm,ҝӏ�Ƽ ��X���"db�G�V~�;���13�3]�F�����>k�G����R��H���Chb,_>�uȄ_�&W�83��2�1�T6A�c��N8���J��²��T���64�/�l1ٿ��G�ǉ<�<WH�!���J��L�ZI-����Q��ş]N}}{��+\�9��#�Q�/"����4ًgbʭ;(���.FV�M�X�O�>���9�۫�@�?����gr1U�^e B�w����:�(m��/�FH��ڍ0���\�*��m`����������+���j^m7'���Pf�lU['Űْ6�f�N���.p�u��f���f?��z�>�Kl^�O��9l�Ǘ{��Du��!i�_���%���!W[��tsL�dA��x�A�d!�Jl�����H=�h3\m�,�������K�X��ԓ|�e��.ˡ--P�8p&3T��s\�4�)H�,x��z�F4{8uo��k�I-\b�zY�n�D�{[(�d�p�MKf@6�,3<U�������"m�YՓ��#��ђCG��) 0��O�����`����*���F	�Cn�]�_x,�W!6��qcy�N֖���v�U���.��8Q��s-�o^�$1Z%XY}�]�5��vR�"��#`�iI�*B?=,�s/63y�΃�WC�L=�@�v�/�2kV]`���2 �c�NvU�����`ҟA�ͺ�?�!�g�R.~��]�B*]�_OVʙֈ�M<:��J���|�@ �h� 5�Gx~���Ek��5���Bf^���<N��+�����S{@�Gn�=��5f�2��K�?9	
(�2�ZH_X���4T'�Uu�V?)��F���,Tjۿ��$������7{���"��G)��M*cX��J�s~��N�e\�۶�����&˗����)<pF�[E��F��1�$4|	[����,S��+�@
#��j�b��[V[R+��껿zv���:��!�lV����73��7��:}}�됖���Lm�9���굂��[��|Z�e,�႞QT���f���$d���I4�ˏ$W���_{{��l)B/(+Q�>�X�B�A�n|}�d�"/
#�wN�է�v��B�qH�� <�
�׋X����^�&��f'8�b��nC�ػo%@h�X�
^��~Y���x�7�n�"I,7k�
�PH�{�?!ҕ�ףʾ=�W�@Ej�"��u�L�}�e�F�s�V���Ao4���8�~�W��#E����,�XJ=v�xE� �ԺYe��l�'t1A7L����>+bQ���h&�r��W�B�Z�mG��1,����y�P ����ځ{YV�7/�<F	��H�+?�9���ݺ�F�_	���p|v6��z�����P��U����xF���܎a�	1��r�fl�!�N��)�p����4�K��_3��,��� �"Z_�jT��iq��ɒX%� ��\9e�GD���f�ǭ�6���E�"���QV�$��wA��H�£�Sd	����}�Nz'�.��f�r���=�-�1R?�����Y'�r��Xmx��G�O�S��3��C��S}an��������y6��{�*k��B*����@�L����O��!%���m�pctVx�w��s'�a_/����Jc�!��-�������p��f��>���1�6Mm7��tHV�5�+�u$%w��u�{Wk4$&�88�?9;����C�4z{(�,�3�c��n�
�c�˄)��Y���`�n|+��\��ۂ�8"�X��~:�G���Of��-��K��ЧLR�!���'�|�⃕��7~0��ǀ�wv�dC�$Wb�)�h�}���/�!��+q�m�e}}$n{N��FRvz?(}{�9�!���G���F��I\3!G]&&Bʉo�!4�,�#�^��g�T���w>���W�:U^���j?��N<����/��gJ &pƞ�V<V]*eW� ����(���o-椛����n��>�T�
���/QW0e�f~��d�=��n��h���F��4�zq����p#��fOI�B����˅Z|��p�(����}�~Ƃ�v�����5��^7��A��|�N��_o���9�Y�J�H�����Q��$�A�@oD�~��w�鍧�-�ڭz&��I=6K"
����N�!$�~�t�g��ێ���l��f_��ݓ��?��z�}�E�I���o��YV2�&8���1g"���F���X�3�]�7���rb�2/�|!!d�;�i4
c�8@w<�u�z4*�ut�����.�ݑ�}���0���s�.�a]uP�mMw��\�\wgۣ|*c���V�D�O��v���/&�]����LXV�(q��$�z���`���L��FI�sv��?��{��]��G��!��+ꊥ��T�D$i��ł1�2����a��4ɉ�K$嗿sHw�<ǾH�@�А��	bD~q���C�y+�3}|b-1�;��ZOSLhZ/6��&�<�g$�y�^(�b�G� P*�W��R���8p��#�Zc�i81q	�����2����9U��aם�v�s��8!|���^$,ny�?�$"1F�q�A5#JI�OփM�PZ�9���А��gۮ���?��t�z#HD�Y{qh���H��Z���b�\�%'>x�Y�1B�X�����,8���0�j(=7�Y��s��X	M�m�g�
"zf����X�^�G5�C5}W���g���y��D�Y�2�x���q��D䆔�;ĕ��7��6�d�?�o��ۈ"�)�Y�� 2)�����d� aڃ%��~AN�+dEu ��	�|���Z�)p#=�OZ
���k�q�:�9��LSY��g]��7?e�h�[Gqj6g~^k�tTslӎ��p����y�����
��^�W��A3�$�%����cN����>�\��I9�D�w���־��p��Z��������Ю�=��g֌cOK��S��o��/\�	{�㥇#o'2@���+nz��,|�R@�,��Mf��49H`��!��g]�/���K���u�J`k���}�W���߽T0F2�]�*�\ٿ!����ّ�)*�M�G��;(���?j�fL�n�!:X��wqLo���.jz>�1�A©3�5Vއ����C��W�h�k�䭦�x�[:��������5n-�|D[�����<c�F�ouCO�bs��}c4� Z �0-��vF=lQ{��W>���le��s��}jYO<XƋ�R`�j��J��r�{�2��'�Q�w�1z;/<�?����Z�Ǐ��ھ��������QB��K[Ϸ��HJ ��2�/����ҝ��;���,/��]-j��u-P&� V��E@)����!b�M�P�aZT�uu\:VB���+�U�˻X:����
X�mM]��ǃ<XL�}MІ5�
�݉���*��<���A�$����&F����,�a��6�O����)��ۍL�.֏x�B�M%tC��c�D�a�<ﰕ����a`dl����n[�K�4�^�m��+}���5�8�<s]�؎iSu���Y+6�\;⯨�,�Em,Q�Y�����=Qst��#}A�=�)�����W��c�W��(Yj�(��ֵw��TB}�x�*����upI�Ah��]�є
�.(� �\��g��I6�?`I	UU�'0H�^�6Y����Q�#9"�Ff;�k552����kN-q�c"fĠ��@��$Z��O?�`�ݭ[�ZL�YU�b��.�juii�dz��ez��P�N�D�>E���.v�c"y�갾��E����T�� �K��k�%�����&{r�ۤ��r0��C�^�)���r�W�����BvYv;��5��+��B�}�Jj8���_8�.~QB	7;�qA��dv��r��&c`�U8���:�^�HS&�6�5m�|��;҆#'�f�9�'*"=AGm�3p�r��*Ӽ���CF����I�dO(ۮ�S��mu�$�H$M+���э��M��])_�qD��>Q%�n��
9\/���Q����<�쒡ZstH��=s=h�t�ʉ֑��>�#-c�݉�����-\!��W�],k�K OF������&��	�)�Rֹ���˿M	��$&���Ⱦ�䋠Y�X�cz����_Ә��Y��Fd�	��C��-�R�\E_�qT�h`����F���������⪖ b�P?�s���0o���^���SJ�1"?F��FVT��
?��R�|!��S��9����Ri���F+�R]��y��͢����*�_x��d����[��"EڽH�ۺ���Q7nc��ڳbt���e{5|{�V��b���*�[C�� �k���(
~��%V�y*��EIIs��#��4ǣ?��DY�Ծ�a�)�/�fN�ѻ�{�+�̛~8_��|s�vv�xی��#Y?�S��X���y���ƙ�)���4o��Cyy뙛��i�	{ka�ቇQ�w�JFY2�L?�^]��Y��6����Q��Չ*>g�ŷ0��I��6�������S~ϖ�띗n��ͯU��O/���	'�[=@E�^�6�F��y�������޼9�����/zk|�P�=��0-<9[�h}�Of ��>䍱ieGJ�Nhy)4��s�j���L�-ȝ�߽L:	���pr�����T(Y���g�HsfO�I���ń{�x"����^U.�h���R�p����+�Q��?	�8����8d5�5Oo�y���(�r��U@�����#����a�5
�n�:���cHJ�З!�/R�G!�k�� 6��q��o�B�^0�6?����ؗ�.��Η�ˠ��S?�+yv%y��܅�z�v����_���I-���?r����U�(���v�H)5�M/�.��8&p�	� ��!��կG@��M��o�+s}�kRaGZ$EK��!�T��v�z����_�Ğ4��#v<�6���V���uqT/"nӛ�Z�:�����Q��
���pe!���.�+ ��Ỉ����t03�#C���
�58Yp��vS~h�M;U	a$��"��1�R]��6���(�4��v<�%cWQ�m��Ó��2$��h����xI{l���O�|�;�e����^o>@<��f��ە��:�jJl�����~6y�T����ǳ�Z��k��̊��%�n	�+"�����e����D���;���gb�n��C~���it�y������>��h����('��T+�SY��SS��=[WL�����~&� H�6'��[yp>}�2�$�,��1J������e���p�fz��k�`�2W�;ەʩe��w��Y���5�����-m-�Z~���x���,��Ii���O��~�(OB�:����.�AgF�i+�S�k�@����E���ׄy���&�
UVa���7TiX��m�I-@e���y���6j�}U@�YE
$o���q�AN��^���=GD�٨�~���1��B&8rjK<��{���w|�A����G�B�ԧ�����~�ʳ�AK��Ǻ�c��S4|�q(:l�N�y(�Go�F�U�s�6k���W��'f��T��TogY0Y	�!�������z�<<��O|v�����q߰3§(ļ,Ȼ9��FG�BE��s��O���sC�ε�Ι�c����f�Ǭ���Ě�j�p��k�~Q������
j��[t>��T#���N=ǭh �vRx�Z�r�����A$,��n� ]��zE��e���~���ѯ��\��J6�Oq.����rZY��6�v[w|�����O\��>Ḱ�� �
z�������g��K2Mu0w9�[`��~㭯8Ҭ�� �3h�?y�\0�@=%Z�a<�dZWYܙ�>e�kI�q�W�M~m�hY!H١z槡������k0Ti���n͉՟��c��(�fG����������jO�v��g�B�5�<|��?D����g��ﳕ��P�\d���y_*؉LC_he�	9�HH=��K>�G�s�@!V&u >L4�}��.`����x��K��B�(J%r���c�7��m�R~	|�<l^k�e�l�a$��1�����h^O�zF3����d��e>AF� ��:ų�B��m����kx�+��mԊ�3��}��\�ο�� c[\H�mm��,E�]��e���/�Z�q�"�ѝ��Ol)���_���U��v1�6G�d����h�������8�������v��D�h��hF��R�v���y=8,�������O�6�L�"�Z�!6����l,�Q%7l��)ނ}E:���0��4l��g�r����*�'&�����C?~0�Q��y�y��}R���ӣ���e-�lg�z�6�[��\���OP%�Z*,w���e�1n�����ކ#�$(� �X2'F�LB[c�ݳF��b�~�5���O�9��m�x��_H2��v_l�H��5_��&���0"����ӝ�ņڠe`=~`��������@Y���?D] ��%� j�
�e��I�_o�X�ے_�\ҼD�-�?��}�0�U%8�E�b5ds`0~U�ӱ�I6[D����&���V�f�c?���!/ ���nx����6�U~߬���GV��o�%�ے,j<�Ӷ��o��Z��6���R�����Q���O;��T��nP��{\�!�Y?�a�O�gD	c�
��@G�rd�8��|2�\�����2�y�kh���cٖg��CnS+q{��tCB� �D��aץ���N���R��xA2?��㰽�(�ݫ�'�N����SA׻pO �t���Ip���C�9!�����W�����%�}��zoߘ�'x�8�w�Pf�#���o�=��+�goy	�/|o<$A�i�I�;r��&+EA ���Һ*hY�E��~GH|����,�!)-I���O�gc}c`Pa������D��5��0���ad�[���������'�u� ����:z�N��a(��<��򺄳� c�a�-g�ן|�U4��铓�z|87��m��_f��ﻏ`
.j����Q�� ����b�8R8������%䆇���/*�Ea�Jxȧd���NYOq.�
�?;n{���L^�8H�Q�Z��B��#�U=����@���A]a��z��)�������'aV�b,dP_�{bX����F���4xcUD)Ѵ�y�3y���僈����k�&��G]���M�K�#r4�-pN&8q�V�V���R!C�m&��4P���ҹ oƱ��+d�W�`;���������I��|)�)��1�O�u��JA��"���T�{@�qVؑ�[Z� y��%����F#�c�T���U_7��ŷ|�J�����N�J=��������Λ��Q�r�7g����F��h� (�:�ڃwd�1��0��>�ѽۼ���yc�$�"l��i��]rן������Bp�CQ�G��@��ߣ(?�m}Lu�+�?D�M���)��h_���	&+�T_�u���m7ժ&/����TROk8˟^(^�h9��h�߁D@^�/a`�a	��w5�خ�f��\�F�F�,�YR�le�x��y����d�gR�h���^6T�tt^=f^]|ɖ�|��x���]���HuP���\�}�`�i�"dz�����"h��짼g4mR�u���n���Y��Y�~��z-=0��.XXʐ�TJ)��s��J�r����z���.Z-g�\�h:�Ɣ����}9:k�<���p������C���W����?7?Mw���+�ڳk_j���9=���*D[��E,�j�����K6�`��BQ��%��*��E{j/�p����a��4L=,���,��I����5(�����1HYi B '~��~V�7�J�=��q��粘�	tL�u!4�4��}��}r�<,.�K
?��gvx� p����e8>�b�*=e��\?Iݾ�t���䫎���I
QP����d	)��Y�m��7���ٽ��>p�Ip�7���|�)ŷ89�w?:��� K���O��?,��5�+�	���Kb/`�Vx�x�M%�:n��i�)��Y�d�,e�i.��E�,'\��um���a������P0�L]�g�I���GY�M{�7/bGL�Zt��k��?��s�@t�
� !��l�īiZ���O�'���i0�)q?�My�O�Ra�P_zN��+3�����6R�H�ay�I �ꁿ�VV��{_Nk�6&^ϊ/N���٤dD�6҄B6�+k�c!�j���Nf;ƬlGjL}�-���O��Ӈ�%v<F����ԈMG�e���/y�%C���YH���먝�,�o�Yˉ��+@G�[�k>��N�����J?�κ�*8�|�m��I���jK��-�x��d�T��y��׽���Xǁ2�ę��8ѳ�Ӱ�<�M*Û�0��6Q!b��Z�/1ၻY�2���k�hA������M� ��Oo��Ih%�r��ܳD����Cc:��*g���2�+���U�
����A��L�3�:*Q6���o�2F�c���8%7�i��i��=yo�񪦶�S>�U����㓸����,�L��n7׳�뮊�$��o �p
��W��g�sT��7�D���$���;n\�9����Gx�q�6�G��հ�(I���&�:��!;iφ�a�Mz6{fS`k���_D��ۙ����F��6ͫ�-���7��Œ)7
S�����~N�vMk��N�7�8o��v���\;�d���m�^��K��,|��%�j[��X4H#W�����-1�UE �=�Z������w�E�N�jڶ�����ʇ����t�9}��;۟�xm�c�H�'-lm�8�;Ah�?Jr���1��n0GDcx�����2��6�rJR�02w����� �A���j�#= .sbY^��i2�Q�/���\���y5v��}�����\��W�YT]��[�󨐏�v���4��U��d3���5��g��B����b������>��2H�;�A6�����i���h�m�<NE�z	����Q���/���Y�!��Q��
����|��ob=�ͬZ�=W˺T,Px%"�%�rV@����'B.}3�O3]y��!��߸@s ���Tvנ���浛瓻64�����L���%:~��!ç}���l�esۖ��HP��m.�����Gnx*�y�Rq�h�7�v��D�����,EY�z��B����g��m��C��_άxS_*��Km� �4�����A��kxH-�i��~[�������S"�t�����dW���4���o�|F�ho�"�[W��v4J��y����?e:�5)`?�gz]��6lY�5{�-�甁9���h�m"pܽ����ثT��̹�^�z�N:;��I��5�FG�\}O��L/����eU�#>8��4�6�m�$p��eh�j-�-�^]��i���$c�m�(�i*
����M.}|y Ǔ�b���xoX�+���������� �w�5�|=?h��,���5N1ÒS���r�A�~}{���N�����E��o�K��d�^�&��ױz]�
���v���V|���q����T��ӇG���Z��xAO�rN�Z(�"T��ʲa��
:�o;�8��`Y�,H�EY�%W{!N�����N�^����ù��cu|L�k��B��MΪ]?@����*�l�X^��"��;�$�ׅH���	����;�E∦���ݹ�#ZD�d �>)&���d~G��E_�D�]d���~���>�|�����p �ku��i��
�N �b�E%>͸2��*�y�2%������2 �6����@Ȓ��\Ճ[�f�1��4�h��u�v�����202yU�����M�1��������D~Q�Yts/��`�~��&�κ�U���FyS�ֳ����J@}c���+|sU@���@�lq-�(�h�^�Lֵ�u�l3�c�d�h)a����59��2��jGk�{��:��Ml³aǷa�C��n`G���ƽ�҂����c�20�a�_�}��m[��ٲ;�5�+�x��/���xZ
*�p`�}<� �5�ɫp@!�j2_Ɔ��rl|E�<s��lP�S|��K��qv��&�̆*�@��G�Pp�R3�>��F�t����e!�cN�[T�f?&�����&�:�/�V%��Y���.ޞ |��c�q��z��c��7}D�E�� �x���������at��7��G��E��� VBt�����8<�K�)�+͈��ڼz�-�q��4���ϋ_W�>������"�n�'{:�ŵ?��C����K�	9��!J� 2��̍ft�b����tݖ\�XN�y��o.� �x�k��0�A���?��vst�|��W�\T��Fk�m���p}.K� )���%���?�yGW�8��A�W|� 2gTH��5N��'�ej��{��W	=����^w��	Y���R���m�5x��������I������RtW�<x�JP�h�9��J��_�82��ʀ5�+9��n���G\u	�z���P���=i;j���y�U	=	2���J�aғ���㪌;6^I�r��l��Ͱ����"Y�wk"��KΕ�����y����oL�&�9�W1�6iY�t���1���UL�C-�ZO�U8Wo? �����NjǏ%����w���=MRaQET�v��X~vp&*#����K��m<�|�,o�|曈�=�Gvs��/�e����NQn�uCN��6)�� ],�V=��JS ��_?*@}+����5��A��t�/��Ng���NҬU	BFM]a3���87�,N��@�Ձ��q���zvU�v88�2;w@k\R�䱻ɛʻ8�^u*����؞Qi��j�%��N�:Y6Ǻ�]�u
��*�~
�we��(�'*fM.Zj��?t���$BK��,��������`�F���NK�{Ւ�_bo�#�QqNҞ;	m����б� C�CxRd;ƽS��еK8iN��߄�D�R��3NX.��������El��}Ԇ_`F=I�>JX�������^&w%s�KiS��t�f��O�T���ѵ�zX���3���ե�I��g
�ſ~��ȏ��D/c�G��J�29�)H_����L�xP����!��H>PG�����<c�f��+��Ӷ|�*��H?���Tx*�	�~�C���v��p��N��,����.w<�t�O���м������MƠ�*��dz����ޣu�s�n�s�=d��%���.��F:zbV��%/e��$F�*�hZ\i{_Fv�����M8Gِ���*�~T�ZrW�L�n���R��Yʛ��}kW�n�̡�檴g�&�S��T�꽙�#��Z�����v�b�G<����|�}�j���u.Sis��=�^��8?O!�)�Y�6���H��U,��u�l�TK���#8']$e�������\���>��{��w��5��jB>%S#^��(B���.}2H�=TO�K@%b�����|]J�?V�	X�8�l����*�7s-�3��	&��(�) �|�_c�1qC�@�Z���wgU���U��+S�E紡*�h�8R��EG�5q�"'S/�'��h%.V�~ �v��.��J�	�7,@��~�=���3O��B��SY#�	����)Csf����!�Q|1V_|��cT��b�����2���■�e�c#�Y
����͕~��F[�	�,aM���Y3G��FD�D��{5�m:���yA�M����sn�|���$x� ٔ@U���d���M�vky�"�"�^AyFM���`���ث��%q�����c˥�r��G�:��r��L�����k/��͓��p��71�(�K�uB��wπ��ޫA����\/mʲ�Z�r���T���"�r��U6F����醲<R�>F���!�^�s�}��d?�l�d.ل��\"�x�mcn��%��	IH��F��JЅ�#��8��`���� �47����7g����j+ %լ{�=�m+B�;����8s�iK�H*fJ���Qw
��֗�'!���������AF4 g�����q@)�]����6?4t�
��m&��!re�d��=�q�
�ӹ����9ׂ�z���d6Bt�����*�	�~)|��Ř(,�l�m�uX��dJ�O�ӹ5 >�d@\�7b����e{� (���7?��.�'&{;i�����v��Ӕ��A�� 5n��KuY�'�M�	��}�z��9�:��$�I�`nv�?��T/��Ĭ:�v�i3�0��/��Q:_9�'����.���\�3����>���r>P4���������ƶ���n��ڎ��I�
�e�֟�A)�n2*��T�Ӥ�4�b�f�P���(�5A�%K��i�@��DS�6��yZ\�-,�V��"�T�9�&�ڃ%���v��i�?���fl��ш�0O�!�_łۉ��C�f�J��N��xVyrѸw�+�_KsA���7����y�4��2�\ꢾ"$d��k��2��+uZ�3D,���U�lB�ESJ��B��#)��U���#��Ŏ��O�
���4�p�ݡ}�_:�� ?pV�\�W:bڦ�4.	߆H��t��UJ�'G!��7��O��Oۇk�$��ϢO�8�d֬�<���"(������ы���s��I��Rsaݸ��0�r����o��M����MTڗ��zߠYնx|&襤o}$��m7ŕPRw�J<��E�98Lo������b��B�8��?@�?�5�3���lԽ>�*�� �>�W���g 0��Jć�"~lM��[�'��L���@�;D�<�������D���?�.��a!�g����u���5+h/zw)���_���ֳK�~�_�o���o�Y���ұ��9�:%u�`�ikuH=ӧ�Ŝ��#-��٠�A��������ŎZ�Z��Y�!��_htz��K�~�y��w^�*��LB��d�#���������o��J�c'T��^p-�g��ݰ��J��<����p�ǔk�x-������|4w���>��E��H|>s#[=;U�M���6s�=@������f���R׶T�|��Y/���.��Bw\��*ʁ��1�j����o��4ۛp�<c�t ��gx�{����"��eOU4g<,�`[�T��U*�:�pS��D�ڽ�y�yu��E��[�WWo����R�� #����k���t�_�?���P��X��LWX�����m/��c�l��h�>C���k��B �Z�X^N��N������]wP�!	}h��N��8{�����P����$Y	�U����+�J�D"~�U���Ի�v�\�z��6�ߺm�z"4c9��5��v%���`��~D;��@NX�3�d�:�t���!���V�^��y`x�=�f'Z����'wk�d�h���d�|����sY���zw�Žn�t>��)��FW��٥���ͽ�u�]�
&���f�S���{\z���8�qג�=&��ƶb�[���3���b/��6�|�i'V�լϝ)��p�NR.���Dį��S�._v�2W�u[����ʵ�(���8H<��	;]�����Z������C���!L���p�ᦕ�v�#>�����q�,�_���s:�Ux���2.ј��[����4t����̛��:��t��4�����������ۣw�����$ő�,�;�D�sOw]=�2ߴX�	�;��0��[-:����X��.���\g_ǩK�F���r�넣̪Z��t/�&>Swt+b��������y��T��ژ��zL��S���ΔM�+w;��+��]���>'h7�yN�0Ъ�#r���O������8]Z��zr������Mva�`��`ҡ" �R�%D@�A�k�6a��` S����" ���ݰ!�Q��>��>�|�O�s�s����9g"V
�LJ��O+��
��f���Tخ�PЎr��U�Z��E�#�0 Ʒ*�m���Q	^3�4��n�=�c����85����QM���)Q�lE6�6��B��Ş�˿%�lPx�b&��g��M�@���/j�Q��Ǒs�L=�{K[*�X;UU�'��"0�^���L}ܻ� ������Y H�!ӤL�o{���OşU�>���r�p����ֺ�P����{�В�w�x�{����
����b-7{���_434�#�U�s�1*32���.%h'�$E2�:��P�zn�Zm[Ps?����^�b��:+V���"���2a:(�����Ϣ+~o�J%�����6V�E;�詫�J�W�4�L�N�7G[yWi��*FW�F.}x%��\�LRG����O�ՙ�J��|���[C!�qS�Z&�q����`�K�j����>�0��/���t�KC#�H�=C��D�Y�A��L��ت����=��C_�w�2҄�F|������o?�9��#�@'LWwc���b3�c�����x�q�c�P�P�g�}��(���6���m�T�4?�ߚ��}���"g00���S�M�hR��%diЅs%)��x��%�)4��L~t��dy+��CIr);U�Q��Jp}B�绿�rKy�'��@(��i���}F�_�0H�m��TN)f̺	/�=AS U��X:c]u����0t�,;�p4�f�����m$͵�G��OmKJ;z,�R�/
��2f��A�>,q�-͟��a�5�s����x��cVw�xC}3�O:6 י�뚆c���0�����4�u��<|\?�G�1g��(/�0/3,S��KS�i
�z�P�&��5���Ĳnu^G9)�(ֲk�D���]���5�Xz��Z�zMn�p�uX��h_��$H�(�_��C���L�PliL<�!����Y�u���Ih�R��(e�f���#��NbF���큕�8���?���V���� ߳K��=2*6�96��!� �ʴ��|PV)ڤ�j�]���F%Pj��O����1hv�$�~̄�ë=�\���~���#a����G��KLz(l_��|��޸q�[Fe�����"vg��Lfc�=��\`��8��>��<�&��],�aN54��������t��H%�q]��B�B,��PY�@ �ni�F���0_�`���&Ŭ���b���0��R�iB��P�t��k`�<��Wc4&�ϧT,��Lhn��>�2�cϾi{�踣�����!S���ȴ�[���V��S��O�A���A�$�ZY�5�Y���I���~T��8�(�k��c��S�r�1��4����Ҥ$��Ӹ=z�8����ӪȓH��1��7t�Ŷ��5bt,�E�1ǒZ��W������o\��d�k�:������{�{!�|K�T���@Z*����(���>�v/�0�//����5Ja�rj.�M��	w>L~���q_��4p���E�>/E�[�e��v��&����L��=��bEϑMj���a��nt���>�H���L��?�B$XQ�r�霝����(Q�TK��f�C�ki/#�����J��~�w�_�b�*2�.ױ���(h�m����5��G/9�����)`/R<ϸ-���������k��h��f�Ŝ�<�،4���d��h7���α��]��02L
V�]��_����>��:'?���]&���Tw7\���$͙0���>:h�w[����lxl��S�Q��QT����@1��]����R�=P����T�j'o�Q��#�H�i#��l~�t��N�5az���ysBQŉ��v��{݉6�x2���|@��s�?�va��<o�e^\�'q��Pa��B���x^���Y�H˧��E�2���!�7���+z�iF՝���q�TS��`��j�4�P�N)�Г�q|����G�^1&��4o9 ŪD7	VI_ˎllQ�Dߝ|��,����o��M� ��u�EJ=�r��&V������<�: ��dy��<�tS��/5j*���we�덛��#�&��uHч>�N�_��X<�^�˕t��Hr	��F��f�5d.\S��;l����~����y��v�.Y;�t�]�g�Q֥\4�v��EF~�ޯB��:|�3\~�_�50s|�UWùW!]y7�T	�Y/���Z�(��jW)`y�J4%�Rh!���v���������ܸ��6pC�"�����ۛ��'g5P�Qy܋oإ�nvm�_�V�uU�d�TUn���(^t�6$_����f��V�Z�&,��9K+��Z��+��,WJ�i"v�e����w������(��>0�f�h���?{�G%�}�"�{�I��5�ܧ��~��U`�,��TU���FNA��S�����n�a6}�\�T�=�S�]h<�3ϡ��(m)�tV���K���( sVb��:˦[Qס�kv��'$�jq�籱X�6�V�r�Mk��I��� �3~���t�A6Hssg���ػ��� {2���咴��r��v��j�'�@��<>��4Y��y;����6��~��̠7-�1�M�xi��tz�.�iVw#ȼl���I�ZZ�̸ӱ�5���@p��i^��E�9E�ި�o�'��M;�_Pm��l��'~�����ʿ1Pu)f��ݾGӛE��;Z�U#�Q��E<]` B��V'��m�"^DR8
ܿB����rm1�$�^>z����k�^����#?�kW�����}SR{�UצoO>Mc���ʆ�K���Ҧ= ��`-�K���M�S� Ƣ¦�_P�Vg��o���Th���:�Ή"=6���pv�9�������]8Qq�`�>���P�_�	u��6�G<������b%��(���f�y%��s��JXE���� ��͠D40'���ѵ�c�M5'(�m����)h����:�c���}H�3I5�e�	!�X�{4�]t���/n/?�)�4g c���S�2���1 #KF��;=d���2s�[��2��&�a{�x |+MSH,�-��܂5��W݋=�&E�]�:�;���2|��t0��e�"~]�k,�A�o���!]�^ �=�2Y���͝=0v��d���x�'�l7�2k��B��*e�"��5����ڱg|��$��y����=��y1t� �ӧ������ű�ĩ}��nEr�*��.�yg�O�]������v�� �}�@�3}������yvmI�������۠F��p]�*��c7�D���<P�0M��������@a�����[�:�<��xX�U��y��+�Ҟ4����=��e7�S`�L��ݨH��1\��;WC�� g��e�n�[J�_q��;
�@WĶ�m�.1��V4�''ιV�P�<�����[(<�'�Q���$-��8�Vk�S���Y:	�5��9������J#�R��R�&͠6!�U���#�H���}b?ϊѦ��zNQ)� J�Bk?%���pr�����Hu�/F��������E#9��j�48�z5nikpg�.�ȴ��_5'/���1~��]���W��|���6�ͼ{<{���P�@n�����Sg��-ç�&�h�3���tN!�[fu~Л�yK����M�"O%�a��~���5�ľ/7�����'������V�'H�emtR�jA ��[�v)��E~>aџ=H�\�[����|p��1>�����u0�t�]5�
�N�z��jr����+b��:s���&�eK��}�&=����z���e�lJ���Fke���b�V��&���
"��6�@j��%�u=�U��X��(�9����?��O���rh�?���O��=��F7k��V|��eE��ˉ�E�	<i*�P'���;g�?2C��>�122&h��[��������`���>Ҳ�Q�
mg@�e��~w��E��Cw��"�����zh2<ג>��&1s���9��}��=Z�p���NցO�[X���+z�ߓ;�'@@�O =�(���ӎ>�/�t���5�J2�|5�L�Yꗨ�3h�-��<!^��0�숡�d�{�sv�z����GEV����+�̰�?��t����6,������/Ts��=}+9U�5��a��眆���	v�I����ِ<ǂ��yNNW/^<aL9hu�k{����=M���O�A6w7<�L��c#ffn����g�۠�?�dBG	���}��	}Hs)<��Chh�ϔ���ͬ���Y��������O{�\�����||��׍�y�����e2�m����D�߸���߸�>s�q�����q�Y�c��/&F��iZ���o�4M���B�2�<;��w׽,�Hi�8�M�z�r�r��j������W��@@5��^�wo	aQ�f�6�F-V��z\��$ׂ�4�_uS�9����oT0��7�5���֮Io[��#�v��_C;����L�!0�k��?��F�^�^�LY��ǡtS�+�j��JE\`�r�s�ȭ��	p�-tր�hq��6���8/��QDRt��]*_���*E������z��{[Jk��9u���y�k�O�%c[i��7P]Q��T���Ly����[�����T��Ȃ�AB�R��n���F.�4x��u�[�oU�ǟy�|&[������O6�~vk7�La�V���,�?G�!N(���s�-�	[w��'�L������Ꙅ���X���,~�f�I4D�%?()x<6����Q���>8���Bf��ho<��݌�U�u�O�����ؗVY�=O��_�9��ӀN���C��_�2)��̬S����u���%Y~������h�h*����M+�\��Kg�Q��͝�=������\������� �G�-R�c/��r\�6'�v��ð<�!Z�~��o�:?粳��U�YHa�aC7��gէ�Ƽ[�����M�1�����CF�O��W쬰uEw*{e�!&HI*���j��t�\����h��EY�����͒��Pr�uS�� E��uY��!�۶	��Y팣*��PD���;`U�1�� ���E����9�N���VA9\	لQU���6w�柩�%5�w��r�P�=�P��lX7W�p8G���F���J	���=�2G�F�O�_�/�n�]��Z5-�*�I�3R���r����Ć26���綍�n6�B3�v�t����؆����՗alBޫ\���u\���0uݴp�.6��a�왠�?jAd0�^��-|\�G�76����n:����� ��ڊKws jyJ�|�x/�9�s*��ԣ�Lq���I�$�ph�-O�H�Ņ�O�(7���K�Wؚ*�k�D�a�@��������K����ذa*V�,x��^1�i��hǖ���x������u�&
E\\?�u��z�-ly���K��B�[~����Ty�)	>쪞�v��sr���n�W"j.��R$��7B�Mɇ���I��+���Q��'�Z���+1�̵��'�r��Kͮ]��>ɂ,Qyf�>Ycc�7�:�9�=�������/T.j�E��>M�t��>o�#hs�М��A�����N��a;�x\�硺+��DG�-	d7��+Q���iA��ß�����}�&|�0RG-�ٮ�_������(���Irݏ�X��Nűq��kS��h\��],�e����?�ݚ9�O��Z�>����k<�}�o$�U�,r�g�Gu�w�w�,���Er�P�i���Be�p�2!�U?b_@�ӝg���E�g���6_���w��"�ȳ�a�4?��w�ij��9ff2�\�T :/��5�OJ�_�=;��i��HL��JUQ�Pj4�C�L�jc���a�h3���˟��IoyKX�'��VG.ض����E���Gkn_���1c,y�H0��ۻ��.sϑ�@q������v�'�-����&"�z�nZ[=��]��^h�]�������7e!.��א`���O���{
��o�5��#r��0*�r%�h!b�˓C�V�p��I�����G^�=����O�����<�yy|kF�g��I٣��q��&?�
��������k�<����}8��x��Q��y����Cz|��5o!�b,�^��#~��Ͳ��M��l��7��6�,��B���z�诮(.|��`���(�u]�"�2oXtY@g�vNQS�@�(|&tO[��.fp���4���YP�T�D���1�w��_��Ӡ�(��N
);/	��@q7-qw���f�ٔ@�� G�k��L���K_M��}3O3��W?�;&?J9 !�p��^�*�+bJ�kF
L$^b/���R*w@��C��q�َ�3�/��Y%�)mw.B	<���l�R|�}��T�SܷH��p`$e�V\C]�S&���;���W?��V9IgG!t�[%�ڗ�����L	`sA \��du5���U� ���f��Nꪠ��P0Ҡ���(d�VCCe��T6%��I2��p�ws2-Z�5�vt�KW!�F��P�oJ��1�ܓ�<n"Pjy�[�5PD�������?qg�Kr!���cOCV��Z#}7v�yy��%u{�uu��u�%���`>�y�fy��g>Z]���H���z�6�LCw�̶��ڇs�J^�W��~��kol��;�^4��.^T)#⼗�����V�͜�`�A־�J@��I��Q�N-�*H��M-�������˻����GV�Mj�!����+d*�Ɣ޻7YV&$��"�ԍ��f*��3��#�������O}�E2�P��;UL���+͠�2	��R��}Mͮ��C[\�t��_N���wg��ʂ��'E���]b��y۠ݻ=k.8�d)f��
v���=V�Q�団��
�{�VĿ�R�����j��l��҇�W�L�qhYfJ��j��[^TU-O���E�����i��>�?6zy�+�EjAB�F;cD�|���>�-t���E���U?+[*~?ĵJ�׉��Ď�{���	��'Q�2���𦠋Q�o��b�[�[ҕRRE����t�+Ԏ��_���tP;I����\/Cx���I��D�A�{RI[i���ZΩQ�#����C�_�y��{�𤸻<<b�q1I?Em�u�g�/G��6�-$ڹ�Ip̸6ڿ/���µA/�y�R%8^��	�~�_4U&
zzB�6��jK	�Y��ܼ���܌�%�]+�(ܠ����
�_׀).~��Xj������MeE^�X�a���k��R�&�2����	�E�^��ic0��]��ܐ�:�tԂ�a����l&Y�-��j�O��
�އW^r4�?���9x�C�F�41'���a���f���&1'�$A�A(p.}�c�|�{�'�b��!%߄�s2M����b�UK���
��1�<;�q�$����庼%����V����/d!Κ��+m:�݅�VG�`��it�+�'���I��2��>ZA\R̋���pSf"����Ŧ/�ݪ�`�8�C>�kfG'�|��De.��N Uf�~���Ϧ%��E���w���%��I���E��z����	��:8�f��7P<b1��_�\����G -������0K���!<[,^R��������x,������Vؑ�l����O�P��z�=���r�=��K
*����k�P�Yk��� ��D_8���Q��e�[�^}�"w��NyY����VY!�al��!>^��~�$֕*pSWy�a߷2^m���͆����_��]��������mY�
��2���y������f����{3Q��kDu��|��P�ŬW��pJb��(p�535f�W�N��F��
�huY(�E��j!�y>�P�a�m�P�����XC)럏�b�Ot1�����6)[��t�ߌ���#�`�YD+�lX˭ުm�KX�IB��2,ܩ<�X����ľ`Q�r�T���2�z��83;��CU>���x6�;�=�6�V^����v��,�� �A7�r�<���F#�.��o3���E�H�J�so׻Ū(C����^�3�;BƋOu���S�{L�Q���A!����
�Fl.��_��N���C��L|_UV[��\���̒]���{o/V��!`�9��{&;�i#����������,�p3y<H7�r�
+���m*sf�)$Z� 3Z�k|�g�dR��U$ݽ,P�\��8?��%\���N`+FV&/����S�3�=٤�{���:�q�n���W�nssa��f�{����̿����N�zog�3"C��d���9��n��g|�?���&�'�W�Vg���OΉ�&���raQGb�
2~�Z�Z��2Q�Y5
�,38X���D��c#8�mI�I;-�t&�jO��SU�}7C��}�W�_��J�;�����=+'�g���oLџ��ڟ��Ć��u��=����R�z���T!���o#�P�>�.�K�}@`Ek���~<�R۹����d�H���ޜ^;��=�;NF7;X��ooil�I &�
A�:���[��0�i7çqC�*\N;�I�l��F�۸�������4�xm�8}�=;n��tU�H��F���P��K��$���w]�זe����V�)�&q�,S���<�0g��v�k��#����#�[�ox	�̗��O��h�gc�L�n� =JT)3��`N�n`e�?�0�C�J���1<lG	����4A��L�3_� z�UCk|�mf��F�C��Adߗ�l�nK�Z{��b+�ϛ���W�b�kK����Jv�mR:��z��,0?��D6e��ec*ٖ�z*��4��������]������?W�q�H�c��I�(�S��<&ç��U�$tG��}m��țP׿������H�/�j��x��#��?�C<��OŖ=+k�Z��dm�ur0�w���袋-�4]��s ��V�1B@�Y���3%��+�6>ab�j�U&jm�������i=S�&!0��,Z^�8ڡ2?����Ć0���l���'~"m|��L��0�������vu�c!N���V~��aƚ�����;�'�=�6�X�"���n�U���ŇEݣ�zx��F_��4��^��];W���l�'�ZP4�KPK�;�ay�="���#�G&�M�]�QƩ���A���2EF�!��>���md;�][�w��{�38�s]Eή��`���`�g�� �.�6ɯf$��*À�2����F5b��0:x�u�N#ㆉ�:�nmҪ3\�BD�1uq�#������W�s�j��꠪[[���q�K}yQ���$��.��X���i����k\��TO*����,������0mm}՞�>�o���J�2�ފ~KaҪ0ߚ4����!�&��"Mж+#�6b}(0�VTr^��F�)ix��E�]��˺��-)*��8��8�˦�辽f��V����F���
ޟ5�	���#4innn�o�g�6���Bܫ5�64�]����?mG$������~�!D�cm�9��N�9)�G�D�l�8�>�\���Oe�wԢ4�^__OS���$aIE�4�>����W�[����D��k��'�Ũ��o͙�Gw�>TTth����񫽟�nRL)��%����o�A�O������ƱQ]�w��k�>���`ؖ2ò�O����Oi��=�On$��������cפ�w��N��{���w��ҐHI��B��Ox� ޹u$�W�16컙�ޚ�ܻ\���؛i�.?R��z7�/O����w�ɾ�˗[��#��4�6��nƛg���R�.W�Z9	"�.�oW�.)�.~�~����U��ӧ���dk�Dg��>�˞-v�&"�\�of��{�YW�a_Ae��4I]��	�H�L|��"⮷\��LK++��jϥ����Kɣ�ie�������v���ĠCU'_��Ș�������n.�9�莢 _�W~B�\�5�rw�2��{y��}����������حsGx�^W;9��R�b�D�r��A_]h���Q_����#Z6i�:Z�>��xh�s�r��Σ�a�
U��?{�L6/�P������:���g�M��E��g��D)�~��{]"V�NK��Z�Nk�7[�9���:�F1�cLݴ~�1`������ȚC�]����gP+��+�>S�c�(.��l��x�&��zƮ'a�����@� ���U�d�]VBf��Mˬ� ��F0�5%�P��?�X��f���I(�p���r�R���'k�%ؕ�!�I��W�@w�,"��ќ�����w%Q�w��[9	'TW��S���!�l -�M�k�[BАc73��ٟ/�Wҧ�w���~`����&j��Җ$��"�(l�}��<�MNNΜ��_l:� '�!K��#L
�۹f�a�5���|�;W��
<���6s��(�sV����̭	��RM���>�q�����E^iC�hc�X�BbK�y�ht��j����X�����Ə�<����R�a'�bY�9�*++�(�`���]�n�ЙE�:����Z�i�g�N8A������X1b�=�zF�YF2b�h��u9A�?�2'<��e�&�!��ܟ��	UZP���� .x0�@���o�4����2�2�߄�b��#��ll ��{���(E�$��'<>ޑ���2; Tȟ���CX��9�N&Z0�yoŠ���XH���|�Bs6f;�'2?��3B�}�S��3�z��ti�&Bܤ���:�WA3�C����	��SB�̾\��S)��l�ȋ_Ϭ�N�~P�6`곥SCd�}xd�0�F�p����וqC6_O�OSD�jj������Hx*�3v�	��/o*��:X�-���z ��}��č  X����5�iuA�2��Hn�Y�Yz Rm�G#k��U�5cSY����rV�98�s;��q����&W�lP��R��̪*L�@���T+l'?�����������,�Ħ+CKZl����!K�J�M�bU<S�^�$��V^�)���
�y�`;�0G����,v� (��ԏw�CB����M�}w�|v��OVJ?9�"V%{��ֶ3�V:�C1H�d�̟��lbG�|+��۵��ʾL��=mݽT�nRή�W�O��6�>�N�!<!�VTՇ�F4��|��x{��7~v��b��Aׇ�R}���Yh�mV�������r���C�R��m�Bd����4 N�2��t����,�&�BB�*]�7��U2"�xmv)BzT�s���������k툷����=5L����e�O�*||����A���ߛ�ɗYhx��ޗ�^��9Y���er� ��0QW�m�F��fAl�!��uε�1��.q�	��� @�д,1��)�d�\1uւ���Aj��N��Y��6"\?�PbV��}���gdޙ�࣒��}��BY�
��Y�M ���*� XD�oq � r���H	b�R*//'��iِ��®�^*w�>��*W�J[��X���,����ͻ')����&���5�r��h��{�����Űe6�Y;J7Y=�������@W��CF��&�c�zzY��ҧ�+��� TkKd�U����u��~r`�)���������:����Wc�w�(KGA��N]�[��������uP_sX�}��NW��_�=����x�ҕ��_�߹D:�������ׯoT:ff��[ooSѲ���F3X��@r^(&�y���G���a._�'�\�r͒������lCCC��.Z��B���W���C�/ �+Z��k�y�,_�/ �Ĉ>V�:g�W�k|l8(���4�s���`���i�V�]��cDl�x�?���n��A�����з�C�|}J���ˀ��d�"""��3��<�t,}�A��H<�,�J|1uƳfE�̈́��߭<����GN�aű6֭Gv�v]����_����T��qtBH�$�}���=)��`�x\-L�����^�8�e�S�C��w�9�����-�����㟼����L�v��x��� A�0>|�Ȳ�c5�r���ƕO�H�(S��o��6�u�f^�!}ma����F��й�s��{8����Kc'k��6w|N���7+��s�Fv���p[����,����e/~� ^�qՐ���:'7H��o�F��$	U:0��C[f2�9{�(�8W����������w)6)ң��8J� ǕWZ�6�ݓ�����#��z���˫�U���^rYMd�˪�.Ğ~l!��5C����g(̄��������=(iN���O�L��t���}��:(C]�����͛�D-2���\��vw��'�Ֆ�EH��d�� ڙ�͜Q@V~��T�����!O��z �F-.2�&����lz��!%�����;�bx�Eߋ�B��o-��F?����.��ս�j��M��~dYU��u�>�
V��ɻ-xr(o�c6��؅���y���Kgr���~�0��{�~Q��d�y��zFa㪕����N^�A�A������0N����^�	��y��A���4l���x����~���PuN`sm��Eg���V}!��#@�}AcE��*����u�����'�����\_� �߷�N��af�Ršдư�v77C�b7�_��;�c��<<<�����ǩ�<��	�u�o�a �]ղ����#��g#�6���/r��TEe��v���>~r������?�%
`aV�]Lgx\����sp��2���p�@�O?"�B�u*ԍ��(nN����R�B��y��s�zQ�ϝ��;�M����DQ�����$=���9�����R��V�/�̲�����CyzE�ϟ�Z�F����;`��u�5 #��N���V�2����j�t�O7���[ic0�Є.�#K|�[K�n��;,s�&����J�[4��6F&�����V�4x��V@�3��D`E�t>]���9Z �5���]C����~]��^�̻	e��-,/�!����7<�T5��1�q�C��Pw�\��$�hJ{CM�+�6�#f�G��H�~H�] P�-|[���.R�M=<ʀi�H�+�}v75������O6 ����Un�����p[�Rd'�>�$k�h��hL�n̰9���;F1Ӟ{/F��7��sdj���#�O\G�y����Z-7ww�B������H����g�^�/��kĽcqa0�����R�ߌE���d@!�{�.���esss�T�Q�����-MMm}����*{�%��<��bb�)h�[w�U�߆�� -�~Rz4~}y|���ੰu�G��.6i~n��۫�nh*eC�Ӟi�L�(f�{y�(?�	q�!M��RYV���A^�͚�͏�'֏U�ͯ�2������&��	�r��v��|4�>��x���%]�&G;�_�lM<��H�ሸ�=v�ϟ?[x2�\�Zdeo��0޻_:���d����e`9���h��y&%ؘ�<����,�'hbع��g�@B �[Z4��'�ؖ���~c�a�p� �_}Cq!!�7o�,����7�fgg���ϵ'�CX�õ;T��z�<Y=E�u�f�x������9�v�w$�eh��k�!��mݻG��kS+rǒ��:���8RJ���Ä�����5�ի��6~�WԢ��EVM����z�Jvv��M����t����:z&Vv���:��J��t�p�>�Ѭu7��v�H�G$����^m�2�� Zd�w�?��r�_��( ���1��e�ei�kk�G��Ⱦ�ۃ�V�u��{���5�ГgΜ�= ���̥?D��ݕ���%C�Q���"���HoH�#z����9Z����**~�Z�1����!���� 
���4��l��SF��W��퉱9�	�Ǣ6�����{qE�>~��(���[W�#�afF��]nE����KyE���PGDF�O·0
+�ϵ�xDn�bH]�հ�-��ND�ō��&	�;w�7�ȸf'�:���ʹj6�h�����c4����mmm��14,��ٙx�H'�������BTDD�wG`����g� j�
�;�x�L.ZQ���\\�mϞ,u,�M��"?��'�t�V8nyh��>@a[@Y7/o��omm�����m4t$'�n�h~6�Wj_��ȴW��G.a}W��(S�yZ
j����7��ؙ��ߊ3�~�s{mZNplhj�ҶX�͑�ݯ<  �������K�E_A��,,���x|��DbP.p)����o	kuH���?���ЕYk��H.y^=VD��^�r,\yե���5[�[]���Tl\�V�p�BB����}3<,�B$���X���0��(q�jY��q�@: �.ǈ:D.--��G%1s� �]ܣt'���'3rs��0�d<qE�H��ً�<=����A˔�4<W�lf!pl��a�0��ǵ[�4�1��!<t�+.�'*��F��n{�Yoo�M0볷�Y%QtJF�������B�6 �:gE��k�8�E��\;��{���smq6�NK6��9���N��^5���>���˟N�t��;-��`�[�ń�,����E��J���ّ����������Ԕy?XF����D4���Y ��Y�_vAA_w����:�ڶ;�
�-�JF!�%'8��e����g�O)�;P���Hȝv�'� ��G���*�O.Lp�Μ=�4mCC�a�wէ��w�qf�!�� R����ˣ��Z�AE\��J�����T�Q�M>'�Z�0H����^�5t;t��O]�0�g+ř�ݕ2��o�B�6�x��2��+��*��L;��nO��Ui�k�[���a.�M��N Ys���F>�7�ࢣ)�#��7M&�@U�]V�o~��礤�I8�����.��[j��66v�y� 	��3H$z&LE[K+!S���;k�&����`��5�1�hA�B�"��
~0��|C���7��#�����֣"�"��"�2�P5����v��	� Q7nj��8 ��H{ 1��5+|�e���y%Cjܔ��x�g*a����s��r�Hdۀ�ɰ�	!��
vȎ�h��1�F
e,ؖ$cVUU�z�+�<��H:������O��o����'�*kL��sɥv�]zd��ࠁaǢ�z�T����_0\���GG�����㴯� � YFn�.3�^u�*_����1���iLL��Ң�������ȭ�5��U���;�?_[�ؐ�]�8)|�������7���MFU�����8L�e�Ú����D�!�x��5OΧ9�|�|
ux��chho0� [*ib�x�"]HQ�c�9�h�0��R (5��K�7�b.�xy���D��tl�K��@F��f��B�����5� ����k{xx|V����HQѡ-V�N-H�j*>>::��Kc��r����Iީ6�����'v��5��(�,�Ҧ��ټ��J�/M�,��Y����)h"׎7�"�
X�}}Z�:-��]`��%SO�Ka�q^M���_޽x¾��ƹ2@7:�6�z�}���+��d ������gM>�g7M�`%ʪ�GJQh(����b\���@������� �k�tq�yc��$<���tt��a����������e���0K��\;�C�aaϿi	��_�,�ߏ&T�����8̑T[~���iY����W�s�wwuu�u�[��k7�̓�-@~����L|��}i�5@.V��7����Ǐߟ������O5QT]}/Wci,��{`)���Ú��p~����g;��NY	Bq�<����z�>��'���������	ۈ� AN�ܢ�����?�[7�kf8���@)�x"���)��)ͯ�>qy�����py ���İTK�Ӏ�;���S��M	�_�Ȟ_�����j���q���1�L0��W��T�5Wz� ��f�g���"No�����_�Va���pǘ�Vtp��Wm
��� �����'o�9�.�o�����4�Y���H�xys�jqN;@G�~}�!R־�qA?�z�#�W��V����.AũdXP\Nhٶ���y��&�.Yx����TE]N�ߦ@��}��κZyX��{���]22�&�eG��Q(}����n�����^�f�����pB����GqS ����b��W��s���d��kX��ӕ�.H�,�~�a���K�wt��&h����/\�մ��}�l���ut���K���j/�l	k�X���1���fG,�;����MU@Z V޴s���0p���"dk��,�	�oh�/�v�_��Ý��A"��sr��h���7A��N�9>���cϼR$[���p�>��w.��z�R�����I�����3���n�KH�f���}��; w����W�D�@��벧����٢O"� �#�4T�Lx8sV�����É=H������ȇ����g.���{��[G�b�O}ɨ���� "�&xW�Z�|���%*}T����3���ǖ��o�ǃ]+�M�^�^a�?�}�}�'�$T����#vYt�xJs�a"��am�{���,^c**�B���:o���٘�_��h �*J���t R9��3e\s%���JN]���V�I�ǶO[-��UW"_�dv��R��}�{�4[0�»�̿s{�j��s'z^]��أ����F��	j&>[}-̗��f��qa�ff7��}�-��� <)~=��>)��%��h�9��UHMP��sj�/Q���:Ƹ�(�r��RWİr��|�����!r���w�L{��ϐ��C��ߕ��oB��� �מ
�����O2,�{ȋ>��r�j3�R�Im������H\�/ـ8=�
��S�$O40,����̉�� �j��	G��<���Cc�IlJ��U�c�\c�/aB����9D�h[���v_�������xٯ+�l�>.`\�����+�kբ>���`����X/��f�F��f�֖����߼��B��,h������9���°G%����y�9��k�7۞��$ɖ΃��\*�M9��oy��=�ϱ�u3s�1k�͔=��J
��~q�k]����GE��=("��Q��/�_�p���|%���J{
��wǈ�YI���P�+����'5!�L>��2+ش���0H�6�'zJ�Hv�42���efb�u� 6����c�â�pQA�CA	II���K��c�ED@����K�`B��AZ��߽���8���Z�zW�}\~L0i!��l�v�^Dt�v+X�ę-���Չptϼ��}���v<%&ygܔܾ	a:�����Mj�!_�����ű���.��Q�n�a/�b(��Jڑ����-Lw��T0�[�-����d���B�	��� �C�XRRM`�O��і�k ���	��g�Hފi�Lt'J�[k�����z��G-}R���\Q�d��H�B��U�2Y~�Mc �⛮<�?�Z=EJ��:���T�FϾ=ظ�,��;x����=_�����A�h]`����*�׹�W'Lp~���`�&���#��j��JRQ�^At�z?�ϳ��r�v ���f�-~�UƼ�����k�
a�.����d��EMtv���:���?�1�o\��//5�Y�ٷ\,���T��U�����T�a݋�Z��|�e�	Vg����̚��u��T���y�D<�� {�5Ȅ.~��R0�pڦ��ɰ��_����¶��)�pU��-:�d��G�7��`Y0��M��*d�������`dˍ+�8]��L�d��/�`p�똦)F����:�D�����u�9���� ��fgw;��N�`�9lY�y���зi�!���{0S�Xd�Y��]�7d]ѣS���p��L��� �Y�ܣB��G������/|
��g�Ye�I����;.�t;/(�n2�~�GiT�r�G��P�5������ wc�����,���>a��*3Y�$E����͌��������nu��ڞ�������Q/�ŗ4�sw3�������n�:�v����7�#E��;κ>��e�8���4���ŲR|y�e�s6���ޔg�R?庞|�c�f͡�gN�ܔ�c�$}���P|C��C�j�U@`E~�)��K��0M��l��\���f��Ν��>�����o=�q����ޚ'j�6�G���7HŗL'~��F�vw~J�R4���p��ЛcV1/b��MAL[�,`�0=�n�"�&}�t9�i>8<�ty��뜚/q�&�eU|f�@ˀ��ɡxG��̟��\���/��M��m�Uttt;X�c�[���B�ҍ���!����7	��-K�V:�Q���g+���;͘3��/�>~1��3k��{e��W�>��g�4�P� S1�kw�`����x��+-+ hB���Ud���Kww��dcN�J��+�|�����z���dRFʓ���mvϿ	q�sFG9��)��a�4��0�ͻeN(��l־��3T�t�ߠQ)�՝Xq��|�阧zbpqJ>��N�Z��OZ���2�DDEK�Po?j��6Л+�3`/�$�C��ni
c&�qV_��G=.s�0����u��v�`4�9��}�a�bj�������Չc�vj���z�ZƝ&�������Ŀ�S83��l+��_x}r���Ҿ#����7��IŢS���c���'�+��^~�u�����#���la�777l�9U�5�i��1v�Vb�V�^����mJWϐ�Aw��U�ڴ���{ �_�[!5�#������$Y�_��$߽\<L_<_�����W�
��a�8:F� b��z.�QvO�����M�����+�O�̎�^����g��݂9��޾=H���3+}k���K���+��C)sM8�T�l���{�M��.[]z�ʔ���뽏�zG�26�Z��a��N��*UDD��w����Zw
e��By����}�#�Dȸ}Ŀ�+l�ϖ7��;%�����G������P �� ����av��$�Cu�/�0b����0�|��G(�y��x&J9���)C��q�ت/污Q���%L��=�S	NZ��<��7̓����qa2�<�k�hښ���a˝^E�q�>X�:�?�|CսU׭oq����va�~���)H���Ӄ^u�T	��m$I0{DT��zlS9T�$�M7?�O�����^fz��
��}�ذR{��-��W� ���e�̩�(e����O�x�I\~���rQ<��:�T*@md��,���k+����UGv�Ͻ�%�����h���'�p'%^��z�20CM�$![��������X�m��/���cꌉ���7��#s��K�X�gSRPR4�Bʄ�?� T�f��<��H�7o�P����������{�_�h��X�}�)I��Z�N���GߏP��������G^���d|�S�,sFv#�C��+L�uP
8^����8Lax�]�du�b�o���G�:͹���@8�w}�Z2"�o<�?�Mu��~�������7�駈a�7A<r�uKO�;A�j����_㜽4V}8�C܏��hs �k�;��P�;D�lnmB���Uz���Ӷ7.W6����c�c�q4_��sf+gO���{�1+KZ��V5��F:��qv�� �{�]��g��ζ4�*9���<��C������b��1���fB��kr��_�/�)j(�nJ�}�E|�ʘ��muN �<N�^L�f$��YK?@-�Hq[X�H�F�,8R���;�~��HN9���BT�e�fw|��ׯc楅76,ŋ�oJc#�_���(o[�h�����ցG�6���#���M�tQ_��3j�@��M��o`3���mB��0�2!�:�$��R�� T�ֽ���Xn��l�����H�䉯4����u�'�n�
Ɔ;�Vpz@��WW�Jf"�5ח##P��zګJľD½���^���Że�r���6,b׽C8̀r����]����Z�7NNf���T����얉X�i�Q�o�U!=��2�l��5������`70c1�Ɓ1�"�wD�?2�~aM�t{ĬuF��p�6�L��j�7ˢu���0>���n�X�)�������<�%���==%��ׯ�|g
�*�_��P��B��8sbi�~���<6�1˗=_srڬ|2��(얞����ͻE���s��V5���Lzd̍�j)ޫ�t+�C_���WY��
Js�[_��������Ӈ��o�a����� �+�(߱���d�h��#�C��;�f���z=Ft���%3,�ɇ͡�*x��!Ld�Z�V����V1d�T��%��aԇ���|wE�/ � �Eػ�U���D������f,�ܛ���d��?�ڨb0	�֫J���#�|p��1�����R!�����?��n�p0;#��;�(�јi�&��T�#mqL�t1����.����o����x��˦Em�� `؂sP<�Oܤ[�����v�3�_�j�D�
�����2��l�����b�
ۢ��9ob9���Ь;>�j�]����쉾��79��W�īI:Sq#I�QK��h���@j�ez0ѷȔ����SP�P�� �k�`�Έ�ϻӢ�A?p9��p�����!1�?�~��"�~o����vw
~�+����$ew<.h�G|�È�����ԘSՍ�����=^��>�wV �Mި�-�Lc�{����[�=d���brO#���ᥲ��u��Y�w8�ޭ�:H̤'�����H�Ww�<0�ǭB�+��z�����=`��' ��^�>�P��������Z��F�L�T�C	�!N	?Ut!�
J �V|��sSp	'��p�殾����������Ɔ��c���]�ۆ41t��k�k�,����"l�U��M[}r�Q�V��kXjTH4�w�uX���yM���?
K��w��%j
c~�h}����7�a���zy�����L�C��2����"��Y�N�S9bA��x$I�L��n�������_�2��nG	�S�ſ5��m��
grKȏ�+� �*m䫩��Mw��g쇚4�]|�ư�W��V�5د��IY��ہ��N�CdNnơ��D���6���ܬ�`^ctx�ӌ�i�F:��y�|E�ʴ{�z�)��P���|PG5oF�8g4����O$�>�J��r%�E�༛mCH ����������/J#��L҆o�E�k�t�c��Yp�޼H%�K��Z���.����;ڂ��u�� ��Ƭ�pfG�Q��M�&,��K�+rU�=I�n�/I���2_��մ�6���Iݑ,+�<S�jqXޟ��h4Z�@�z�T-3��~��z�]DP��"Z���v`������:ң�y�$���R�oO'�t%�ڏ�!�;kf"u5E��]�qe�!b�[�~���E�W`p��}1�ťD0�	f.��<k�`��j���m��%�v�˧�j��w��27:���eԋH�3d��шJ����[�$���^6��O�3���>'�"S�`����xxw)�.<-���N<tmI'n�@6�(N�ް�U����=��+q���#(4�t�U]�.X�%4�<ls��N�|h��B������9=�N2}�J��h-�E�j� P(w����ct�|�:��r}��s2�2��md܃�*7�9�٘��G��!&UB�&c>����:�G�|�<��u���;�����س7��\!�~�N�����c��!Z��}>s�]��oJ�}аz3����&x��͌ ����ܢ�)d&7��-�Mo���*��[�J,���PcВ�������b�Qݬ�b��4����	��$�t�?��Ш�ٽ��K�׿�y#M(��Y_͠�t�iPs����,��9�*�/O#��k��(��إ��0��v�'�eZt��:}��^����(R��2�b��&�=�G9�EC�_j|a���g��z)������g��\!� �y��-#-�R�kV��a5)t4�Iva�����3c���EY_Ϣ�E����M��f+�����!+�Ih|�G���W���v�l��!�,RAO����oN��8O�Z�����I+8%_@ic�gn���DQ"c,�m,�x"�Dh"Ez����'M:��{��D!����m2�� ��b)�4D�ƫ{S��N]�H���'fΐ�Є���t�ޑ�n�v���*�g��eV0�A�~$?[9AEa(��A=�5���Tux`��Up!��e��Nh�����U��E؏��ĬTd#�gj*+��x<�i��yv�U�`&�.-w���/����&�����+&D�r�SO�\��*�����/j7"ݾ�n|}�����4r���� �^��|l�=q4����_<=H�nL�fAA�\||��P~uaha�:�;���PS�E2���x1;�CK}e�5����S|�uoCI�o�ϣ�h2�A�p���8єX�G
W�U��U�h�l��T���(��o��6I_V��5�:Z��z4�X�~�iG��<u��|�8��MU�0B�5v�Q�p�;�����I
��(��CD
������`�>��5 1=_��2*�<]=Q�^�iN�t��J#r�B�v�tJM���C����#5$�?�rj�-,���.|��$�I�R!�8+@�?3|��NX2�n��{fG�������%׏��{�,S������Ͽ�6���G�;����hg4W7��1A�Zd_��˙�9j	R��G>��P�q�k�\��L�:���q|H�V=�����M/U� ��81>ZUKN�e�s-�N�!eG�iq�9�{�;7�l��Gs�/.ޣ�
�wgΎ��꥛}�������6�[�h
|ErMqf�:�<�/�u��8� �K�U�4�1��R)ð<\���������2��]/	{ ����$G�hp���74*�d��~���Tl�˜���$(gb����Y�4�b1l�.�� ]�;�^�r#�ۛ��)��R�ϷV������16A|�`|���C]V
�]K&�Q�
��qJ�(:�tSh�7�)x>��t��+�&L���c�!X¹M��`�
�/��lf(��I��:~0�Eeb���q��A����|َu�2�q}:�A�S��[o�ͪ/_*�!�t��ɼ�����P`L+&ox?/5�
���b�f��|U��"�ħd"��Y��W����Nye5b˄�������a��0*�Р/%*$Ѳ��X�W�Th��TZ�xrx����l^��b�	=�r�����Y-��Z�xi�-�l����b_�'������%�VP69&�uJ�D���m[*wf�vU�2p�v�D1�N.J��� ٿ��@�b/��o�mm��N�j������Սu4�-�W��=lw�7���أ������E��yt�T{��v��T
D���R�e��dTXÌïga�/� +_��zeH�'V-3V �^װ�oY�v���9)�M�~!�-|�N�H�����p*�8:����R������N\�c,��=r�P�5Cg�ۄ=�>�?,��<b@�� e��Hp��?D�]�������xg<?[D��B�A�R�dNEzXC�;���u��{�$����I���O{#������L�i�I�g]7�% * �ga	g3���>�g���ѹ'.�h��E=	���J�񓪔����z{���2^�@��r�Y�EdN.�8�)�[j9&�p~6Azi�ٟ������|���@��`��	�����59z�M�l'�|R�N_��)3?�nw�@���
��bj��[B ?y�o�0��R��Uw	Z��e]��J�P8.�����&$��f��ɣ�K\ X�H��/�?	̢�aR }��ւx��̑�Ң�
�:�d~�2����uw�؍����jM���ǯ��h^�ϛ���ə?%u*b����k�+���`�0/<@լ�>ei���F�Q�v����dH6��.@N%H��ɼ��DX�����7-������<�>\K���'Yc)��	���׫\�Vٓ��T;3�p�;���'�~�0'ҦqPƟ7�$$�b��+���l�u7c
|�#��AE���g�C�'#k$PQ�����헝\#�feO2d��q��u�m4��.��������v,�C���K̜���K��,9a9K�~p�Z�7���S��$�B��۩�����%���R����(~9���o��3�E��5?�.��u�_��>G}��q����W�9ɖ���&>~==��8_F�*�R@���7�Ʒ��2�������-�۽N\�PT.����pv|3���y	���a���F!�%u2��� 0�	���c��.z]������
�d�}\�M�<\�YP�j�/a0j���b��$pz�f�<f]��wNNg,��0ۘ9hv�����j���zkŭ�7�j�10׳>%����<`1Yx3���Hd_���� �f�P���w/�̽�q��9�}����m|ʵ9�r� ݰ}�#u4�x#����9����p�7��Wv��N��c۹�3ot;�����H����w��. �@J��+���ѻENf":W0j�g9����K6����ηL�u��ۆ>� ��s�^��
��%��Wǈ�@Y��^��n�|P�H�lD{��[����Ȼ���`=$6l�H�˘��K�Ԥ�(Rn��n>���V(d���	b�˳�.	��#=��j�7@J@s���%�Eu`u�3�97=����}���@wTTe=�W,�����*E����C����R��M�𺔗>6n�&G�S�{�jʒ���+B�?�@�REj����_�X/�@��?78��H����6(��a��r"���m3l���)xŘ"�x�{�i�:��sÖ"�h^x�<Z�Hҥ�J�>ۏ��&6"��<�����F�T�����Y3-o����aX�Xנ�7ȳ�E���[�!P��]�8�ք��VO�}�y�~�����i:��9��p�v�H���(A�r���X|��-e��������^f��*3���b�K�w~�R���n|}���W������Ne㓇��������m��H�V�`�]�b�:֥�K�7`zO����ᡦ~nY�vS"�'/VR��gF�^�b���4�*9w�G)�!:7Hc�ݮԱ=uHE��T�miaz��������L?%� `k222ԓ���d~dI�MC���X��zE��i�Y�
/8��6pP�nDJ��P�'�ܩe^�l�K��x)�UG�!��֢~�Pf��[ �C]��l�!w�w��pm����ϫ����Z�p�J�t�����XX�-4�1N4�e���h��f�"v��n۝��['I���=�?8���2�.��C�?�|׆+I�Vw�f>�|EM���m[�}����!���{�>�ȧ��'��K�F��F��o��cX�X��7�3���lrP8͏_w(I6uo
~X�sN��
�Z0���L�?W�0�X���2P�si��/�=�\*����_���g�-̝ʴ��Ld]� {"{��MuG���CM-��@����)���-w�a�Lk�X��t�%�8rՏ��߂a���,gRcAO����p���4ief�~7J�g���v�v�:	�d�	`48����e���'�6H�Pz鄮�kun�M�v�H2~at}<Z)�� ���d�^ :�f[�g��W}�UXR�{�Բ8L�_#"2��b'��w�	�5���|���4aՉ[�C��JXҕ=�����n��e?�,��?a4��Q M�5��c9Gk��m��Z7q{�_E���r���OXoW2�ş��xKoM�N�Q,29e�𐺩����;'QS/����[ki�LI��a��cOM����"U�0���,�F�P���W:ŝY���2.�n���Ӟz3�[8C���H��@�ϛ.L��\ի�^N�*9,O�an�,om}z�h����g���ɾ��R(�9���n� �H�烪)|@�!|]j�Y*a����������ަ ()ϊ���/+���{�<��*.U4��8�|?ތ�Fڔ����e���1>�yָ�wZ����o��N��^��+{wc�p����u6\��~�y���Jҹ�wr���f�5����ZO|4����A�Ԙo�()+w���/5�F����Y�����E�/ARL���7�P)^����|_܎j��!Z�W ��;�:�E�Y������be��&�[��Ŭ� v�*���p�{��WƔ)��/�t���q��b�_��C=
��ߤ8�uDf��rk�&l����vz6mUԿZk����zGy����L�fg��U�hk�q{� �c�(�_~�U"��R)��[�Enj�`�_;Z}V��$��>�}]�y�֨��lV������� El��0i�e�A��-���G�K���v�M�|��+C�_\�A�2%���d�������YΨ��m^3i��\��8����t*��)$�tP���Lz�mq{z}�1p��0J8L�����{�k���qfW��M3D�M��`�wpq6$zzzԓ�� Sʹ��OQ9_����<6W�_>�I���u�=Ԝ	����p=E����Z��k��Dd����܂��'���i٫���3e��z�Y���x�X� ࣷ���M�VI�������S�Ӛk$�� ���]=%���O��Rs��{�E�F�/�~��j7*��\��8��Uq}=�~joY���n�*<z��#���-Ʃ����cW�5S���Rm?�>V��ӧM�[+�T��U�
��pz�<o����;DD���/I?�o����pv~��*�d�.n
B���M�?�=�ث��
`���Y�Ǌ���F'��������@��?O%�K��5B��L���T���h�F��u���YE\��&�g�񢗌�������V�at���m�ve׸�� wڟ����^%��"FK���� S���n�Exw�3}#r�i�+�ߣ[ۥ7���˜& m_��L�N(5����"B�i�b	С����� .��ç�TA�oV�=���J���$Se$f�ϵz�#=�cif�n_�(��.��ģ�\`��,�$� ���}"�Y�'��Y1R[_��$��R&A:Y����V�=+��+�����s�����S;
���/��Sr�}��}�k>��3�|�O8���I<�W�v�2�w� ?i}����Q~33Ύ�Yqs��&��`L�e�xg�_�Ɯ���Ǐ}�)�r��W�o�Ǳ����2zƳx��������[bp�Ȫ+����x-�/�.� Z�ń��w����-�3��v9���Lō]�����(tm�[Ϫ��X���d�/�^AmV�0k�K�?G��ud;�Z/��q�T�k8��!�����BppX����`�S�G������3?[- ��N�HI�[�d�UN)��e�Um�OD�%��Y�j��W��σ/�W��,\�����ɟ����H�!܌ΔQ��K5!&��iU����E�4�{�Ͽ������F�FIc@�u�b�D��T"���Swj��^@�*8Ik(pp�y��?7)X�0]���^f�L�e�G�@�M���+**0�$�(���6���m��n<����TBW� [i���!c���P�22�A�]�&��1_����m��V�@S��w�&��ޣ�t��NY?]�5��;�-:)�r�J7����
7b��c(�����doyh���ygR�2@�IC��T�P�;�-Sh���s�y�0�CM�[����DL�1����q؛m���v;O��2����-C�OR���� �y�:��|�eHJd��Ѿ���3+t�#��� t9,�����T�F�S*:���Ɵ��{u��+c�3��X_M���q-<����؝	�Kk�C0�EG���PS�ʞ�d~��\� L���L��V=$um,�����/o�)��h3��a�ʷM�2�F��լ-�,�;rLI;��GWL[�����F�6$�MU�-��N��"W�w(
�^n���i� �׿�M݈ ͙���в-����n��h!d
xoJʭ�����̾�V_��@]�MU����f�*X����o�I��R��5IJI�G����'�.�'b�|�� ���E��=����."�4����za�Es�xĕ�ǿ|&�/ ����h"�k"��X<
䲊Z�����ARKف�S7���e�[A�-�mB8RSQ��|f-$�!I�,vr���-�3"t#P)�r'}	W�Ж�^�s����cϞ��J�ޱ1�w�K.Ҡ��W���GØ%�*��~�Psc�;���S�I��7\SRY%�۝&:cGo�ǣ���*#)���M��������d� s��G.oz'��r�'�x�H �����~�q9�xg�;�{��wJ�:��mi�
Xr5�K�����6�u��~���W���w�8eOvg!�/S%�����|�뢡g�CCC�Ldΐ�J�� �$Uc�h���)�IG!M;���d3b7��ޕ�4ꁣ̯��:���ݔga�&fp��*>H�k6�d�[��l�^�~��q ��=ɼ�>�:õLX�M�������;I�N�Z��Q2�p��I���]�r�"���wK����LC�>��ՙ��'7St|���9[��U����NQeU������5�DH�`����Tu�g�Uљ͕7k������޷n�tD.'O��/��-���+R���˷�6��/L�[��}���`'�^% �����];�Η~<�O��C��	���:�Iß�x7$�w(����S�ː�[Lt\ry;��rT��"v��|���)��o���S��+����U��`B������6�"��|y��V:�"7�	�w���E@��[�UTn�~����e��$��"J$����چ/fi����P�7�D���BYț���k)����Y�w�Qa)�h��{ts7�B62�8kZ-{ ������q����O��)�-F��)��]*�)�"�
=/��~�m��6�=>J����S�ȝ$�ﵟ��>;�.c. �2l����Wg���Nȭ�2�L�X,��cf+�N��>2�1J��#l�q�������c��b�h挕�����z(aސ���z1f]~UsRy��æ�ED��_�T��2�v���h>��ʟҺ�ugu����1�6�7o8I���f�Bv�&��s�s���`�ՙ�D��Ga�m)4� �����#B]xhIs��᳣�Ē�A������QF��aO:/|R���h��.���bn;�?�9�����DA�[ZL�euu0QO�}}�'/��)R�ji2�~���=p�d7�a��;��m�P�,%1�NX����XJ�bTA�ɻ:Jr'�g^�T��Z����Z�e�mK����`e3s�]����i*Je�n�N�f�Bq�c�A�켸u�qRjy�c3�_!Kܺ~� �Q�-�6�oj||��/f��МS��Ϝ��+}Ɍ��!v�6��K��*�T�p%��e_T���)B���R���s���$����墋4:�f}������n��/L�Ǘ��4�i��n4�`��2ձ�O�C��&@]���1�9le��bkkK�1�+�Vy �JJ�l���ˉn�$���co[�w�y�T���[����b�&������1v�7�Xj~�a�3�X>>��6�������Q�l^:�?Թ�a�
��׾���;�KS���OL���UO
�k���ԟF��MV�n̢i"�k3��W���߸wZWL�5��M��ͩ,.��^�3s��~��=ҝV�k]VX�/�������WH��ݎ궀WȀ����~���Dz@��U�^5:� z��-��=xq�S�)M]�r��&�+K� v��d啽���cR�	�x�V���*�� Q�X�o�\�o�ᦈ䤊����HNR��|�7�p��1��A�W�Ԗ���-�i�q5RG�mT�me/i���z#J*qZ�6�eٕ��#�
@9Vb2UR�R �Z�L��Oμ[��\i5N~�������T*���E��zd��>&� 9ϧQ xb�WSk��aC�S�$��@���%9��$9O=Q�:��0�AVo��Q�5e�$�z#�4�7Y�܏CR%[�x� ���G���I�'.(�!B���,�^�b4�{'y(B<0$F�,cX�$%=��kb�=2��#������R��mXB�&��y^���K������I�,�d@|���O��1���UeV�v���B�6��n_�+k��&NXM��1��N���T"�P)����<����3v�no�Sp��,A��������'��.!�G-B�555%�?��$Yt�o��L`c GSqOܩm��S�-�tF���IxИ���-�_�g��J�X@f�̷�9���8���pN�upf8[9�{3��5�w<��t҆�٢N&�,��jHsĹa��J���1�8��I�k����YsHQ_ϔNX���N��*�%�o������r ad�d�!|��Q�p���؋�~͙�Fk2W54������+� �a^rl�I�������X�P`@��	��m�績�B���k̋q�>iw�=ig��Mx�F�l���,�-�����X�������</���c(�*=�w�B���V.�(]	΄y����r�>�0���r�D���̈́�/8����2;���Pk��V:t��`�#��5-�������O��=���#�xfe~ҧ"��a�����J}K=�*r����0��3[�������+��1���*̏�.�.T&#����EUز�N��+��rpp� ҟt�����$�	�@�\�II:e�P�C'�Sd&yBzۭ�΍��2[���FL !���C�������&�j���-t>��]�R�Jw��ʋ{oi�r���ʟf50�W�M�YOA�`���OeGй��[^~��GU<P �E���u���-�QW�U���}�(+��4�߶���-�H`��c�h����}2�%Sx�ppP��wQhW�o`�Ii.�����f�)+�7�i�����'	��&Lat�J�紥C	��L�Ez�WJ���æ���Z<��������o ��T�m��qmY��*'mM�ԏ:�]+^��v�.b��7-��@<��H9�9�8�"�0�S�|�ס����h%�"�;�fz�<�C�@�m��w�3���U�l��{Q�?��Gm���_���!�3$sA`�CK��	����5��J���=+�IX��������|�ᓴ��2�ˋ\Nz��C4�{n�x|�����ø�{�T���&��R-�C,ePc��EE���;#t��Y07蘯��H�SM�6H���Z��'���Yc�?~��vw|�ː ~�[q�*��淵}���R����$_�N�$?�Ec�е ���<���r����V�3v��0�X���;�r��H���m4i)G�B���P�Ǚ�t�ny��|}��1F����1K��|�y���|S����&N����\����AZ�3���������4!���1:���v�o��2ǌ!��M��ScYͶ!
H�2�AB������ZH����I����epP��S�N1�:�^��/��&�.ڃ����7��>�qP�>��uq���:z���;ɌO�u�)x���C����E�� vp�!0S�������������z��(oGhՃ4�VC��ܷ2 ����y&���9N�P��<�s��\9pՕ�������g�_{);`s��ڷ��G�lzsƱ�kW�)��>V5�:4qF��v�8+�B|SLA+<�g���t����)B%���#�O	O����D,�8�a
o8Kf���쁦��iI%ھ�I�G\�YI���}��	W���E=�F��RE�Y,�z�z
���D��^�;��a�mB�f0{��6�l^
׸gc����;�z���1.����&|j�P��M"��JȠ��B�Q���]��]�X#�N�P�쨒՛N�XSc3k�%>%!�̋��*��{��sƉV�N��S紸�ay��G�6̟�z�����F\�G��ݶ�`&�.�j�Bq�_��iU�b�ٷt�Ȝ������j���v{������r���R<�\�����G��m{ӯ=B���d٥�k�m`�"�	��h�5������[���l�Aa�K�򃦅��Q�ʨ(��篞OUm3���Q�a�udE�9c���a$� ���@�K�
P}B��w����RՃ�J*;�V��/��M_7[}C�����'�m R��J{ 9㺮�u
/W&�.j9y��zu�N��d-�/v�U��#+}f����A���S6n:�I.��{M43Uc�B��c̘'a����|8��1k}�+��^���q�������lP���Ycj%�t����H�|�ѡ�'%?�3ir�y<���#۲���W��5i�O���	�xO��Ꟈ����d_�\P9@���E��@����<��mK��EY2|�P��p��]�
KB6��)��VJ�x[�dXQ����ї�����^�G~#jR��q�nl|��^���YE�\>@�z�)z?��on�;[a�Tg�n�׫��[(��|�mq6���>���;cƬ���p�J1堰��U���s�Z�}�O��� S�7����|���Ld��݈�����KPU1�(c�}x �	v���Q�����P�q�\����6�ӣ<�y����$��	�i��ЃE?嫯tehb����;<e}�{s�v�;�\��'Y��~����]�6%�Y��ދ�p:���))/TdͿ}���(�dU��.��
����x��:���nQ2��5�1PE�L�ή0.��u�j�[='M�g�L���� a��:�^O�$-���� �Z���bQ�w�3{����|i�R�\��殺�l�o,-��w�]�mg���KצS/���/?vx�oN��$\�j�x/W�zaRɻ�K4���Ѓ��~Ҁ �ZI#��[ ��/u$�{=[9Ranj��)�Fս
�s�˧���� ���k�7c��qӭ�+	���\�;cظ�軒�+[ޠ�C������i%}�����k���Y0I����	C�QLϱ���6v�N��Cê�!���hگ���8n'�|τc}M��a�Bb���˩�j|�Y���DI���J���v�S�1�	P��$h��Н�{������/�FU��;����g�ff�2���q��H5�.Ս��P�-ҟp%�KVi�%lN�X�͠�>��G:�e�UQ���4=�d,z*
?�/2�j:�}��u�n: �@���&���Ⱦ�Y쾣�N�1}4jl��9������^���VL7R��s9�V7u|�K�ԱGIq7���M��o�w�z����e�O������Λ[���i���@4���:Ik��Z�j}nFS�)�D�D�����Tm+/�#�֜F@f��iN�T�>�	=��!y�v�;�����pq�)���<V�C}����Z�En���ޗ��,�"�!�+F��(�&6C��G��N�}�8C�N�d6Gb�a��-�����$L���w>	��"�s�RD��msy9��yG����e7 R�`l�_�Y S�j��v����[�ӿ��_�|�G&x������@|��S_IC�z��:��|Z�-b�	r)���o$ p�eΔ/���9о�;,#X;)#@���#ɬ9��T[�\�2H��d��6��oŞ;E2�<^j@�1�s]�m�m�/�.�ڀL�7�tTZ�.2_�c��ioOO�9CX�����4�����z�$���tUd�_���)vB����v�Ah,��oR�#�a�YQT��O�U��2~�1�#�9�?�[k�j��j����� �>ї�����^�������B�������Rgҿ�6��>��FBN��%��������?��LR7mi��|�޻6����qc��xĤ�d��N���?Be�c�!�C��sW�����V�BW�NA�S_�S3`�.,�o�P���-#e�N!(&⭌���ﳪ!�����)�I�plCGUS�a��1�,X�=���H%\P��J~�sw>�k	1s��5�g�_8(����������YL��r�z\��$o����wk����x;���ҩ��ɝ�S"Qt��B����J�N����h�:���y��q�Z��nt�
�I
p����6���3�3��Rq�R������~�E����i��6<��O����)���숎"�¸6Nfje�*w׆�o�
�������q��v�����s�S`����4����&x�������{Å�P1h�%��D�:D:�F:Q$��c@����n���o�����k�b13g�����y����	P�#=`�Ɂ���D6Q�۹��w�z�F<�{�?��*WE f>�ҹ��Qۼ�D�f^�}u�H�g2��3�K��l��w�KH�}�}c!��� ��y�zޓ�-��D��O�{���u���v���}JG���R~^aup���O���uՕZsEU�؆"�#6��b��o�Oha2�=�(�o�C���F�=K_{�knI��@� tc�u�b�a!�̡M�v��j�;/�?�m$��|��0T�������j������9ݫh��q�U��Hi~��u+׾�j�t#���v�~v���Q鵌���=��6�'}��~��W5h�#x�~�ޡ�[X����oVM�n��z��*˪�g��[$z�B2����u�^wU�N�'���*�e�@l�	!�?��J�|x�A����@����թ�ї��eKB�)rX��<�{8�8"7�/� �
O�r����]5�����w���[��y5fi�q��h��q�bu��ջ�P�r^��M1[<w��>>�����>�S�/ ���/��?muCK��ǿ�z��y�q<��V���_u9��U�b�R8hJ�w�I�YSkf�C����cJ��h�y5���)��u�����=O���;�.ͥ5BS0uFp7:I۹qE6����P���^��o�5U����0��V��q���Bg�q�2�kbA-�f&jy�?���O�}_b��U�a�%��'6(��W��e�����.=N��_���n���8nLi�tz���/_=9L�D����#l4�a�N|�O���D���=���u�>&�HSWD�JT~�X���a`�IV�y���AJ;j��t�O�=tG:���m.뭍Ķx%�������Oc�78o� Smss9Sr=%ཹ[u�� ���%g��y�ԙt��s��Me�z�+M��~� ?/��t��t~���+`$IEo�ڃwP��fp��'��R3ݯ%qbo�ZZX���}���\M��#�P h�I.�eq-���?��~�hbL�e���6�ݳ}d�%��Z�E9��{�ܝb�KVQ��̩�j��M�k�ۺP;�����wrK��:d��ٲ��4���8�:4��.H��$��{{s=[��KTO(��G���g�_w��g�9_�u��<h�0+�ve��`sW���\6���Q�Gυ�����_�ka�{ȼ'9��µ:TV+�ڂ���\挠��������'�2�!4	'R1�w�*��kz_΃���N+�8g*�z�xΖ�繫�N�7��cO�,��R���,��$��N��Ma:��X�r�3bv��|�v�!� ?��C��6��\�N��L��7�{$��]�(T�S�_����H��g�w.~��C�h=g7�G*?�<C��U�禲���L3K��:X�ߺ�q�/���+=�|}EV�3�y"��mo��0��vn� v�vN��[��ea��Ç
1t�2$	=���^3+Ͻ/!�c�Z=��)����{cǏ:<hƛ�9E�NH�h�u��"���qyd��:5�1Kp��n�4��u-.���os�~��'��jQ���H�@��c��V�"Yk��v{�^r�xK�y$Σ]A �{3Df���l�&����TO�^*.��n�v���>,`��w���љ5W?����j�"��\���lv��s�d�t�ٴ`R��6��g	/"������J^�qr3boDD�z�^�?�N݊��h>��~�u*tȱ S���^J)�����-!�@�x��<���	�]joi7ň����nr�������ٗ<�+�t럤"nl=|]� ���;)����F�ۑ�A���ȉ�I��Jb�v����a��B%�x������~(US���e����i�F������2����#	uA	��Z`��V�a�G)[!��X����q��.N;H�?hF0(�z�x&����>2�
Br���c��E^��wb�]7��hc>Rpf}��-�##��qi���Ѱ���LH֭
��7�'���7��4��#W~�������**+w�bi�ܺ��1{ָ�^���˙yO䪋2/OV����b�Ύ'V��	��	�|�lw�X�M}��Xȟ"��j�S�j�p���0�� �4�u�?�z�����#$��9����nG%�P0z�����k�*��G$!�l���.�g�d�%F>,�h�����G�8���9�܃ёV���I{�/�����:e��+T"�2@�%Q�u�s����6K�h=B�^�����b
�8��j��l���"C�R}]�WHk��P��}�7	�U�T!h�X��"��^�83�[��G���ZFn ���^�]��l�a�;.����uU����Z/a������0�/3����6z��#��_zWaw��sۃ#t��N^�jX%,�C��;�$���4�M��<k%C�P�Zl�â놉��b/wz��nK��'�wٝ 7X�����ׄBS�!�=����+�~]�h��:����Ƴdj���R;�~���uu���ou�%'"E��������S�r��!��\z*uc͓�Jtc	Ϻ�tQE��>����4Z�z=�����~�
1�T|hx
-���4�Qdddm&���r����W��p���4DP��OT��k/2{dتm�%$@��g˖}ڽOoSc��e�t
Q�c���f�ɂ��^�YMZ-�@���h˝���* Þ�_j@�cn���"��W@�=�h~�@9���r'����M������0�|�������蛷F!Č>A7�,_H��t�2r~m�&�5����1�"�LBtEB���g���J]�[=?)}oe�F��ƵA_�c��S�Pe��;f�g�Jb�RV�����`��V�k_�	�b�m��s��a��� �e\��}�׾?�(n���N����S&皌����Dx.F����"���Ԙ��<�4�~��� ��Ɔ%	�����2��8��w��T	�8h[�2G<6
��)���_����;K��J����uz����9�0$��[�J.����5�aSz�k��Q�2PP,ad�?�dۓ�$�]7k6���v���D�����ޞ>�5�e����,V��-f���xIQ`s�З#uc�5_]�3�l���� ~Ծһ>b��=­��A`��t��F@7�$9�L�K�{6=�/|%s����.<&#��f�ws�<��/��n�~l6H�H�%��<jߘ���b��/$F��k:��~mE��n�X��=_���Q,e�0��)�U7���N"W����W>xܭ�X���=���433�w�r*	�#�ۮb+_�ܙNɘ+��^��=��N����c��o�����
��]�}�������S���]�-�d�፼��rʅ^��|}��Ӈ{�CX0�y���K����E�3�Mα7���P}�kPr�u|��{#���O3��0�qny����}���CIT��׫�_#R!&s?��`�Ų���x&�e�2������q�F�SI�
���/��Bd}�����ĸ~zb�:O��Zh�쉙�LL2�FL&)�7��ӄI-,,����T��΍����;M��L�����G-z���Y��Ɣ=������x�|O`R�WX��D�$�`�$i��'j��&&&.1���jͱ�cs�?���2�YKu��J�d*����<���/�����������t8��Dd���x_�LLmp���9�ٚn�~pQ�p͜2����J@h��v߮)wݔ�����CS8�d�2k��� w���-�7%2(FDG�"�Gd��=��%��T�g~���}�!j��A�&��UNZ��B���d�>;����_�	��j�'%?}�S��}�T��������ǐ �yF�����ƌ�ĀoZ}:N����D��Q=�[.����q�y	ON�r a�\�=�PVQy���������5����7��m��<z�����%�~L�ðVcĽ�i��Q_�"�E�~Vt4����ks��[~T[-�@���M������e%U�| '?A!;"Bl��A"��ߋbUK�Yތ�����%�����?}y?	�;7�G&af	�p+T^��_�XZo>������́_|^��۷%S�AE�Mi�+��ݚ�S^�.��Ræ�!��.��5�~U6È��M�B�R����@�4�W���3��B���~Wʹ����sr�z�'&���{]����g��,�z��K7qu�<���1_���B���72鈨'�������ǯ�?&f�P\<�\|I����(	�8SI��|Ua��Ic��Os�EyY�*��]�(��ؒ4�J���į��+��14Q�� w�S�/\0ZE���QX��YFł����Q_�B�#0>�b����b�o�35c��+�͢9T����S;�������ġ,/��G����T��X���n��֘M�������eLbgl�R����U1�S���ʩ�� YTq�*�[�HO�ߞ$�Xg{���B�t)�q㟂����Q�������������o�d}�آ4�L���F�Ǌ<x"�-��:�6M�`��,��W�|Ҵ������-E�JG���n5�'u��ӕ�	{)�틣:>���I&��΅���3���v&ՇD��0f���iNQ��p�U�do,�J5"5z��҇�>��`��	�ٲv�}_��	�̂�|f��������O��؀�_���#6.�]T6�q�ґ��Jvr��6����KqR3�2��V�i�	�??�H`qZ�M����?�kg���%&n�¢����UUեI����<�e�jg���w:��;̢t�ጷ�7&*�F��uYAA�Τ�ed@��֨˴�F�c�;a�`�4A 	�ݓ����44L��wX#v�0�f�SW������Q��� �����U�r%l�����o�FQ!�}:䈕u�^�6���"��P�.1<<`k�+e��#�<�|�S΄勩�/_Rrr�P_:���{ƫQ4�$N��6�Nܘu�+����f\&�V��� ��T݆�R��SU���#5�ts1葉��́���8U$%�P�����O�o
j�����ݗ{Ll/eB�͉���z�d���
����-bjjV�N�tj*��r�>�G	�h���Hy����I�"���s�SݽV�b!RZ�9�����\/'����	���'<�~J���{މ?�����KWA�I��߯�~�<�����ǪYL���H�I�JfZ�d=^˪)[��(�f����P��_�K�C#H(���W�+�ʙS�|m�bA���ۺ�<��
H�K^q�V��+)��q����(��\$VV$�:�?+�y̖�߫-i�L�w�݌-�������Z���|,X���o{G�����X)����d�jG������>��E�^Bu555�&�+�%�RJ#���g}�&�R4��?�)Fŉ�l���Ulm����WX��<����b���f�=���!�:����E޻��/4�
Uq�׍�����î�)"*0,�m����0Z7���v��'��	�$�f�@ �M���nd�
u���ۖR���b�����eo�hE�ⵃߤkOM,,r;c��	�8�I|���x��"��v�fE�>Pj:׍ONF�xi�ꑇaV�d�H�:k���%��6Q�U��!�z�hj��1f��_g��4�2ng#T8��K�i^�7,7������m��V�z� p������<�)�I;�.��s{;A�%_���LV�E����n�A͚n�׾����v�����Լ������h�I��O�o�YTH�TO���"ؠi� �jGp�f�W��<����ն�y�$��֟ g��2�T%���$�G��Åq�ل
jAF�$<޶�>�>�>�[p�v��\��B��$�#�j�`"��e �ݱ�O�'�-"��/��X�PB���蕬��v~�P��>G5��u��h�3e��<����X�vl�������c0�)�������]]��Ϸ����E�b�n��n�r�7??=bfg'lw�5���KJ�����׺|����_Me��Қ[��PU��7:���st'�����Q��Ҳ����tr�]>pD��u��l�>��zF-���j9¥'��T�(����r��'�P�^w�O�)�'N��l-�T2�]�ǝ�ҦL$p�q6�t�{;���T�0�if�5���u�G>�ǏR|
�j��VL&��j�\��9���d��"+�?��{����!�h���~%���U�V�g�r���yE2�su����"
���������ܹ19�6��,�)���%�;jF�>т���I��5ihi�V;.Y��YX��V.�����Gl/�x}L��E<��(-Ws-�k]{�M%S���]�Å��������ӑ����$\e����8R�����l��s���W�h�,<���7��j�x��ng�tPr.�>==��KC�+: �JR��o�i���[\t|r���\����OB����Xܞ�	����3��g��1w��i�s&.�s�l��Xt���)�z�B.�K,��B�+��]�˰�(�����@]�u�(��kW�����'�`u�u/�Cd,��1�+����ڶ��q85�q�k��M{�䫨E���y���)�/�s�h�����UWW�O;�'�^��K��a_	�}uk�u�n�u�:^�Mr6���1Ԕ����@B�G2�z��ݮׯ�2� ��Sj�c�~j޲����Vͽ
A���CT+#�v���y v�G��v�N����H��59g�ԧ�d�p��ob�Aܓ��l3£zYs�r���h������87lL���m �h�׺Q��Cd����v��hm3m�띯M�>�����v%	鐑5��1�hVz�n�B��z�gX�<Q!�����;��P�ƭ�aA`��EW��O߲j��	cdB�]�z]|���I�����V��1ޡ�μ..`��s����>>q��K���)ŗH1Z����8��T��Wo��'���� -��z|���To�]�>��4u=n��	/-�C���5�ݤ�G�q;Z�e ����H"�H;�a���jb n����S�J*�bl�>&�
��u?�J�EYl����>L�}9�۪��h'%`ԇ���c`���!�#m �"���գ��׹u*����.3g4��v�K����U�@B����#_���uA̯u]�H騣,��%�B
-�݉�����6��c��>�'�VV�~��� ���2���P�懰���A��넒�t�њ���*5�\˰���$����|,_�Y��Ÿ�dף���!F6
w��� ~u����S+���d���W�L�%����N(�8r��8�.���m�O���no1��rw�+��&�F_�2�p��(�k�4AУ�p6l+uv�zF6�P�е�Yu"��2�Ь!p���4�������S��d�"�c�����u�������~ϫƏ�J����5��Ӽ1�TH�R�#�����j=��9�q�=���¶G�ȵE�WL�~i��=ަ�i!��dzҎ�.�W���cЬz�b�[;}�%%�e���CPQ��4$�
p�O�>ql��*+��v~��  ���n��?'�~4=-��=��ܝ:U
��Ws��-Q26o�A|��)�_y�~����4�⊿s��$�gړ�n�2.����@x�q|k�B׬�ۏ��}�g�����<�[(7�Q]�)(N��BݥH���y��C�xGk-�XӮ8���7ZÀ�iwEJ^�2k/��;q���n5 ��'�������rx��V���=���(��is��U����0��Pi�#��0ř�MAQ�㪫�6�B�̏����k��?��y�Z���=O�
�as��m��W#,��_A�n�ϫ��4�'N
34ŏ #o���b����ڋb!{4��_����m��Y3�;���q� 7�a�ڝ�6�}Eʅ�	���ڛh1��@��wvw�c	�e���x����=s���c���U]�0�����GS����@�ά{���7���4��e��x��^���X�}oY�n�������D��������|�ͪ�+s�k��/��|� J��<n�{K���1��Y��>���k�(�� j�"e�1�/���Nv֛\�	}U>�.</��%�&.�~�l�kb$V/���v��h�%�`^�h���Z����o�^������d��	��E���͑0�>�� �7:R�9H��naϹދ����4�N�Z�����q;:���W'�ή8���8ʟ^Ss�7\!I�b�|"/'穳��Naȍ�g�v�+ӻ�u�k}��Ž
YȖ��jM������>)�ՇZ5W}B���J��"��h�~W�:;�A�w��c�~���<�\��sӗNݕ��E�ۧ$�����|WVE1��lwb&�n�3�a�JĦz��6T@���U+u�ϱ�c׵�?�}�bc����'����z��H���U�+��fa�=��/�)��ĭ+tq�����rQ�4��˘kT� ��u�������q�2�@��j�F.�+B�ޟ,%{�\�������������,xJ.w���%�N<��*�t�l�S�e�*�k66F^n?+_�"�@���u$�c�;��K��
�7V'^
����x�E�S�{��'=�H�|mH�0qU͂�Jm�I�Uߞ XDO��0b�ᗡw��<�>q�f1�W�nW����c?���ۘ�_�1"'����D�rD*a�i�ŷ��ULQ�Gix��o$v�p�1�0s�6��.3AJ5�)��g�P�N4�5�{����Y���9�8곔>`���_����`ƭ�}%������A��!���w� A�ѹ� ��?a�Hzs�`�5����mZBw���u��_�jOG��kx�N�lΘ��d��V����J���j�䌌lŏ��N`q�8�d��F rÀ�u��}�V�u��P�윗{��Pe����v氩L�}�����S&ߺ)M��
�;[�hf?��VY2}|�G����f��Ft��u��Rx�G���t�/��p;���7gB^?U��5@�_�`ZE�É�Vk�[C-��� B�!��[��9D�NV)��a�i��l;�a�߯�����H	<�J�km4aRvg����7������/ۈ~�G���C�s�Xߝ�9J�?����?jPv�����?��y��UMd�Z�^u�)"��7]�%��:��xK/.�P%:���2E��
�;�nS���V#֬3U�M��F����j��jY����^�}}$<_����In�}�(�̴�Gk��%%%��J�[	X�uf��_��	&{�|b�������&R��YRd��m����i�g!���3��w%4^�s>��T$b)�ڙ��*������� zC]�A6.�H��aʇ�DT'��=}���R\G��O�l��g�P.�f�>
`+<_�2���`�!��b�V�{=&�D����~������6��sԍ��[Ă����A�V��b���e�m�"!�m�B*�^�2�N0f�Xv1�pA�kf^�զe�mZcsV�`���v�IB�\n{��˽sAƅX|�
B[�8��aw���Ԗ3c���饰��@�����,i�o�W�!��V4�[��M�ͺ�<�J[8�����?�ϝF�P��ΰ-5��JMWf��cu�R���"����{�j��5%�n���x����t�P�ꌚ`��es�F����$?�g�!���{�N ��,jչ���gS�V5!G���/EmF怠|he;�GNFŜ��u�c���J��Go�}J�ꎷ�7��7R#���%��U2�%*�*�Ro�{=yN�^+[�g��*��Od,I��(Y���F;�'��{v��'BR����*����ʱx��c��|�'y�@��=�y0��q�&jʶ+�W�}�䍧؋-��u�m]>YXh�io{KT\\X���qg������°���b%�_�Sܖ�L�Y�[���;l�9v�G�"0���ܶ�ϡv�G���_���I�h4V��M!�fs�/΅\ �?�}O��M��vu�1�j��i�����n�)55�����m�����b�e�[�����pY�3�m5� dߝ9��L��ͭ�>QypTE�
����c��#�V��:��͛-�i}��_������;�U�l�ޖ)3��[�,�U��B:�k=��|�lt�!�#ÃGU��΁ 6��Qd��+�!'kl8X;nu������#ϑ�/��R��m����=SV͒�?I��Ѫ?CZ��I;�Z�(����("��&j����#4��D��Ϝ��AG1 �a1\� �R�·��ΐ��@#��>[=�fMxm7�]���V�`RC����@Z���ð���:������y��Ѽnaa2��!+'��WF��[ �YL׺
O��a�0����+�
����g�׵m�iw���}���#e�]I)>n�F�#��t�SA��E��[��nl���Uhf�E�R���]�Y�K&�C܃�t,�?i� ��|���c���#&f�~�+7���=��ۿ ��>����k�t�����t��1YMLL��.���	|PMH��${���90	kc��[���1]#�){S��� �T]l;�47.ddg[��m�ij��a���޶t��P?d0�P8{���"o{OO�!+GK�p�Xci��t�DΫ��qPO&,�}033spyA�g�!�6�����M����uu��1�jZ&k�݉u�yg�Is� ĕ�R��Wn�/���Yw9��{�K{Vt�y7��i��j��>����S�܁��$>1�;��<��~[`7��a0�6������k,����TX����v�^1Ѯh��.�c�~�!B;��;V���ح�K����ݬ$h����);�	d/�_uwv�Y�KD��R�J�jk[��iRvY�Zuu����RT��j�rD`�v����_��a������Z��m_�-�j�A��F��XA���f\�Lj+U��N�X�N�u�u�Vms�)�I�a�x ��K����g����U�Ɇ��6ʥpy8��| �]h��:f��}복L����t���h�֗�Xmg��{*+�]�?�͟ogwZ���Wv�Q�ڡ���5�x�"]�l�x�r�]��""�\���b��Z�Kc�xQ�>�z4���}LÀ���m8+j72�vv�|�%�;b�G��ɜW�e�@�Q;��x�}���6���PyЬ�V�/O?�o{�}w�32�Pp֫"�3��_�^�i�I�}h+$X�)"5�����|fְ����:aYu���<�=�]���rַ	D"4��*���s��{:��D6�VD�q�ߜ���I	,c�|��X<7^%}B�݌~�оfc�o���J��L٘2ˡ<�E>�Ӫ;O4S>�2���n_�=����R=q�dザޖ?�ǃ��7Gև��X�H�擹ϧ���`)�]�fs��#���d��7����Τ]/E�~�w6�}���Hp�"&�*{�&n���U�7���,XV)}$����ۂ8Yt�:۵�9z(����?8���z��~�$-��k6�a�0ʎfՁ
���X6����M�wI���]�R��D�R�W�����ITQG�|W|��� bc�Үv;�[�
:r�g7��%�@�ocZ����3q��?�M�GX��w�wcZ�~R�0�n�R��O�T��\3�&��Iy"^��^2��wݹ���$�?��>>���p��r�⣣�y���q�v�/t�={��y/�����U�A�"��׋U�@I�jY�B�x�����]�U�(�us	Q1��������BLz�vQ��m"�ǔ��!��2��}� Ҏ��ͽ/��ՃIHVꏢ��U㥭�l(]�b�>�`G9����PS5�V\�U[�Aw�ȾR�դ|�l��~ΙZw�`��纠��n�g�F5�8�	=l����6|f6?a>R·��Q���g<�,@�l��"\T��!kl�yV�P� ԋ��k�5A�r�8���6��m-�hl����oT�DEG���	�0Ob�?���j���n2��ٛ�D���X��SQp�~

*s?��Y�8�`��x�ⲉċo�o�	�&D&ю��]�e1M�V�x�e���6Z�����v�l
[4��S�,�	l����������`�����n��j6��P:9��Do�?��{O(���ZT����h���S�j��i��<lDk��d�[�	�AF���i�3���N���6)�MO���9��\�bJ\���,�:�#&��Z}�v}�v�X'��1YW�2X��L}ݼndx]��iIX�.5 �;��#C^�*�5�TYZO���n��Z#:neA�Ѳn*^VU�pȀ������̌�D&nr���=�L"n=p��̾����>듛�y��%s�۸?�G�����B�>{�;�DN���`���iO�S�Fؚ���� )��{��c��nK99��
�̦rջ�@P�G�I+�h@
�z~,iC��T���1y�L>��(����9�չ�Պ��z��54H�#<8iq;x��޶u�<�狻8�S�2+c�֫y�1��W={���7�'��n�0��A\����~^EP侭{3�w�(P!y\�2����P�����n}�U���+N�{�}5+Y�klW����2�u+Q�}x�&����Qw��ٜ��;������;S���!!C��I��P������}��`�o��TU��k@��_d���>�;��Up�*Ga�n�q��T�3�m��*q<���|ox�m��� 0mʺ�/F)~k�`J@
��%�L6{�yk��u����X�d�O�[�	/��5���<<��
��_�#"Ҥ�>z��aˆ�����z.���ʗ/)��\�:7�l\�ׯӲ�bŪ���C(󑼊�nT6 �)J���C�e;�a�|���i�˳�w�)[|���S=���Y;�q;sݗ	W�G:!/{IV�ҏ?��<u_%�A*�վ�@pY�/IIE d�<~��,EZVv`0W5��Wc��F�2�>105'.� �u(��ϣ�t���$���5PNϻi|*o�ݭ���і���l���ߜU2:W4�:�LMvo:S��_���E�57����?���P��M���y_��ooo@1߸5L���Nܮ;oZ~�׻aX�����lW�
��'�M�h��\���������pa�l�\\tQ�Kn5�ˈ�,`Ȏ�!���ޗ�HHI1��������$FCz�*�Y��4�k�k�φ�߉��U���|<�|�v9���<�
����֎��,D�Hs�t�G&�ل��)������.��gk�c���O����^��R[ߦ�(s�9���2� o���Ƭܯf����6�l�eQ�=�ieN=��4cccn�K �X ���$!��$w|J�2���/���JԭF��FT�2#oIKM=�|�e����o���7��kQ�[w��7��?��%!����ǅn�F"FfR���$��sWdT�9�#������I�Ո���Y���*X���/�Źa���VCyQY
�y�?��ڣ���`�m+5��oyV#Eq\���A��B����5���4�:���UQ\ ��d����V��������t�xU�ƾ�t�����d�W��3)�*�Q7�r�Vk��}E�#��t�Z�R�ja4B�����[1�>(�a�#= U�B��m�O�����OA H����&�g��`�{���
�o�2)���	/�/>�H-����:��������n~�
ܹ�J�����8/�۶�5;��-* 3Y����0��2��@��Q���[δɎ���t�\\#x�9�U�qS��P�M�J���{�a�OK�K�/� ��jeee��]���XN0��ֿ�ܧ���2�a=0UT�w��R��E�����꫅]מ-������G���nM�|6M2��e?j����f�N���b�l���O�b��$����N�1�&��4�V4��D0��)~n��ԩ��R�i�R$s6Ai`>�ZQ@H硦檦��Kx��DD��^^���fc�
���:N=B�/��m��$~eq����w8=���`N�k�Ϡ�yKK=d�WG*���'O�Kk��Cβo��G%ŧ�P�D�A���d������o7�ф�t��7� =�<��w	(����4��ǲ���%��u�M���gǛ%�y6_�&,aD47V�~�J�C�>x��E?f)&�+�9��f���rv���v�Q�x�Bph�0}� ����IB�{���Ķ�25�������=�,8�(������-�����ݛd����h{�$_b�Ӳ��s�4*
.?4_�A��~���w�;��QuQ]���ܯ�Sl��X;E�T�ׁ�ϙ�m�#�lر��5_U�0�:ԁd}��u��`Q�O!!�1lz�M�~�{�py;��8A������E@`b����0L@Z���+/�㱘���|r���h��3i��!>�Ob���p��%Q�J��Ȩ��IH�X���~�<���g��	r|�<�k�0-��,�����r��Q>�p�t�>5m����s�"N (P�C]M9J��{��OVl��<�0#�Jҋg°X��z�V�?����˭�ߴ��
�\�`��?���'�)9��z��jC��5��fp�(����V�:�xĠ �$�xJ4��j&̅G�_b�tУ5<�?>K$֩i�5��v~���*�{*���`�{�~mvuz�KaӠ�4���6/c~�oPQAJA?TƁ�2VN���Y�n�^��@���ݡm�L�f0R��ZW�����|>F� S`�V��QfU�&�Y�`���H(i��ܧ	��tu���{���W�免2���mh�,Z���5u����O�D��i����&,}MS/;xi#[хκ��(�<JBV�y13R��û�`��Wנ��/�˓�6�͒=M�_
҄�����+7���~�b�ɢQ q���\V�O֧�&  ��;���N�k�|�s'�>uh�t�c
fe�t#b�$y���8|AO�(�UR�֭ڠ oI-p�5�ΎR��p���o�K���w	/?�����A�|M��}'x�0��D��:��:�]�]���ݝJ=,�m��
�X`6W�)� �M��^_��x�M<�����"�[?jΏрJW���zaqq�p{�M~6�Ǣ}�s#�;_l
��)V�7z�MJi�c�"��C2�j�5���z�^��ZWȵ[W&���:<�>�ޥ�i��f��k6HdaR-��3�d���H��(#m��q/:��s�.Vq�Z�y�߉��Ⱦ�FX��������5�yZ�H8�HMZ��BZ[0 ���hˍ�j�w[)`@����3g�Y�k�ي�`R��DD��_��3�n���j�+F���2���I�S.6���d�u*G���f7t]b�p\c���|}PS�����A�,�n����B�{3�/*���?���k-��q�Z���j�U]?�O�^1ꖬ����� $^��T���k�����wu����3Y]_�H9�e�ʭ۸��d$p"�e>�ƍj����MX8WG���AІ��`��y?�_��ɉ����
��1<d�y�BGI��-��7�=��L��W \%
���'�_��HT�zK|ށ"{�8�3?����7Gm��BΨ[���MyTL��,�����3DiW{:
���=$[7y䈱���uv�ܘHtU�4���q�ٟ�C�T����x-qIMɨ{���;�A�Q��\9A;Rܥ�+�jH�QOQ#�n�g���/�7���gi��g\�'�Zz��ӏ��F�P�G����������~bE�T1c6;}�����+�OF��͈Ř�P�����@8Q����o�پ�n�ٯ�aX�������~�d���ĆYu���G�b�v�F0Q��9�����B�]��跇P��Q�,��Y�A���
����]g��lbꚦ>/|�phRzE���]�0���R�)wϊ�s��a�����0��#�	Oe�����J���r���-��Z��K���?�;2�E�(�J�p�(����y}����zFޭ�\جR��T�!/���)?b��w�!���q##ɶ��1 #hf����X���y1�=9�+��\y{{�%�=�ΘY��Jf^QQ�6����V�j]�<���f����	�P�͡���hK�aŪ[)�!�N�������G�:����Uߓ_�3MPx���a����EE� \ґ����Z� �U�v˺�"�*��xU���	-;�ɨ�1��#R�="O�7��b/��2�� L~��S�!�;�?C��}m;7J-�g���~����z !��۷%s#k3��bj>�Ҥު+��Ĭ���^5�\qʓ
�9>F#��Mj�~Ar������灹f�2�L���� ���_���fH��P蘒���J"�5V����-�����Ȗ!��Rg&G��YNj��������\\.?��d>��qڕ��`F)���[�g�h�,���I��>{�^���̓<�/ I�;%���--/?$N(��J��WD����v~K���fƭ'T���E�v0��^I_�m�/�l�סQ%o����õ��j��F�>]P�f�T���z�	^��S}�oSR�X��] �7FPե����^�2$�޸��(�ïL���˘�;pXxaq�@�3$��5x��_찯���3��\�|��e�r����?����{!MWV�T����9��_�v���@_�#2 .���'a������qF&'�I�~�'##�@�،�i����v�e�z�3�T�9�U���,�����q-J@�.��h�7�47�u%�
 6�L����g������Ua�2�k�o���ԏ���4�ew`1R�B�k��D���r���O�Uh	�-b5R9]�V��8����k4�f��>������ݸq*A #�����{�*ƿ>o�������Q��Θ4��=�C�q�Z�m�.A�y���;U��dde�!�2Z�#򈃃c/��TL�⨇��Ҫ=�E�x�E��������ｙ�x�z-���]�����1�*o�%.B��Eކ���V�X������b
ܶ0�D~���J������޵���-�� OA����zP�[J�ْ���U��s>�t\j5Ť>��Q�NgP��C��oN�KJJ(� �v����) 0l���(Xqw�+�cG��:����D������qhhD'�.�����WL��	��M�%�.JA�n������:7L?��ᆱL^D����/��h�$^��ݍ��;������5MLM�99U�)yY��i�1l�"������Or���?�~�A(>Y�L^�:�2�Nȅ����C7��1�PQ����("R �:�tKǐ��t#��]H# 
H3����- ��C:t�������k�֕����g�O�g�3a��5��$ tA���K�:bS=�,(`i<������UX�+����B��yԒ�\�,�+��Z���RB��{�:[��8r��k��Ltӓ�fЉws���~ܽ5+�w����.G�"��
���S`���=����!,��������wɱ!�c�lf��%�lO���]"����,,�!/��ňoLUۥ��'�iK�ٵaxg��P�ܸL��II�BɅ�����^J�v$��6xl"�BR�1f�\��;�T�9�����{�P��t-�Ẳ����u@L��N��R�����������$Qي�m" z>��ꨴ_z����yj[<\�d&|���c�ewA�.��4�����]OM-�*��)�}�E۩@ǰ{��>~��0��zq[}+H�jzW/��K�mciz�H�>/OX����B����.�Q|�՟�{����2�h��Bh���̄M���%5�l3���Vϙ������e-��#((l{�cΛ��:�?�,8�  �Y���E.8�A-���y�D�%K���:r�q��	�8k�>�p~�A|�}_!���u��C쪧{2 X��}@-�@K۞=q�"����*�l�����z��
��'G�$����XXX�|>V�×��4HQx����g�]����/��xq`61��4zc��0P�&ffV=ь�w�'̧+r/�(��A��k���݇�2��e�5;Eiw�J�N|p_^�@^u-��q��ٟՔdx�J��_�)��Zj�>� vsPV�����,���c`{��
�x@�OR�׻1���z��ey���#eeepl��e\oP�g�l����f�~��oKQ�Q\�����~{>z:���c�B6x�
f��3{B0y��h�B�x�%w��&p[���]������m�?Zmg���u�-
�wHG*����NH�8������	�&���:�A�s�/c���SuJ�[������5��ߢ�f
^���Dؘ[�IĀC�?�n���x�'�β-�جI+m��x�l���Z���Ar�����b}odt4i���ܛ���Nd[���x��$p��8�yX���0�+S1�Ǹ��Q��p�����v�ux�������++��	�A3Jk�	�,5r���s���[g�нS_�TY�V�unt:ڹ��F&���UC9�i\b�jט�uc�Cs��t'�h���t����d�>e%W�U�
mf�����`�9K��4�\i��x����� H�M����&��mN�M'��x�V_��p�y�Ri�ꨨ����X�Y,�_{���B�j�����yp�@�q�U������'|�Oh;�oU軘��ٚ���|�!���<��3H��c���
˷{<c1|Q.��k>$�Q~��fW�(����-�c;;�ң���������k�֫�f ��2��@����:���0��fi'��8i������-0K��w�>���
�pWI�<�-9H���l>I��T�ǻ�^Ui�6��.Ͻ�{$g�G)۫b��%�����Md~�����Ұ�.���,�ZMG �k�]n��[Ol�#�\�r X��r����,d1r0�~1=("g0�^ޔJ�nF�E1��ݺ�ׁ,*�S������#�k1G���1(��wF���UXO�Dcu�'��">�2����@>�/�%F�P��у���
��8�hߕa����{�~1��YGiۅ������s	dOdO\(����K�݃<������ۘr��=(����1�q��@�2˙��<��j��yV?�.A�>���c���	����#��R@�ׯ���$�%��֞���i��D�M�e<c ��W��s)�kڐ;��3<j�7o�B�hwTr�h(������5y��?��%���Xs^��;*�qY��UH�x~�shh�;9����/����?�zl [lэ?����ibb��2�8�� ��z��M�`��}\�O3����?+j�O\�z�g�C�_���JPPHJe�H��Z�뉇�I���I,�@�*y���R�j`�H#�+�+f)��5޸a��'�@x������+*�{'jNWq��Ӽ}`w�L�3�-:�=�R߾�����U[�4(`�� #����c�v����~�H@}۶d&m���U�H�պ"�ۢD,�W?����W��dv�ݙ��5�>�����W�"�u����5Re���� ���WFj/�D�X)���GY��8�Yj$�;q��g������A]����V�L�r���t�����j�������3"�o�w��{�t��҈QF�K�G��ܰ�QZ�֖���S��5����$�Ѭ�80�7�\��?uڞ� ���'�F����ð�����匭&E��Z�1�9o{�~Qz�w��C�7@;i��xo(�v1�`������S��\O?a��4z\��4���T7�K�	���Ϫ=�����"�K��o�V�#�8���i�O�Ԛ�EGiR=��!!P�]���~y��X�	����?�ʴl��?�}1Co6[q�z¨�&���aD�:�C���B��ɱ�PĸC�T�'��p9��Cl��%5��(O�Fh̑�=D��C��|	
��9:����۰�����ez���H�ד��ڵ���*�B�F�YjȯX�c�k"�WBJ$U�������'6M����?����b�aQ{������`
���A��X�N3r��,��(�����m��$�id6Y���T&{��l��AF�`#���e�F\�R#{ňu�='�\&:X�@y������A�~�����o����$j��R99z��hh C�����I�u�gh��B+�c��}*{8�&������6&�$�I@1[OU�C�an� f~�e)��%��G�����6����}z�T�	f��k�ғ���CFg�Q~.)���.peM�3C����x"vll�l�O�巃A�=�_��~M(]usë\5�No���ڭ?�7����p��˜<���$Ә��_}�E�N[L���Q��V���ӳ���5D�,=�Q��+t�,�� �)�Լ�v�p��*�ӫ�`��ZS��Q9rvC_0hn��ԩ᭱�@@��Y`-�U�7Fٶמ��^�I�c�����k�o�W˪��Og@-��fu�]j��F#03շ�R�����:n+�Nx�Z���<�r7��f��`�u�w<�SJ�_������/xrB���@�����G̤�!w�%�z1D&2ƒ����a������:�n㑷wIbu�fh��nx�-��U�7��D���\�ނ	���?�y|��K>��
%{�5a�O�)mi���>�,dlluf���ǃ�6hc��?�Ŷ��*��43H��V�<Q�*�*��N���Ux���|�?m�5�j�*���&�Tvy�GTX~b6ʪ�wu�s������Y�oףM���o�E!Z��:�:�*k�����sX ��1o�`���9��k��gK���~�#��ՓG���+_��'�?�]�p%rb���� OF��Fr@F� �

����Aaj��'��~>.�a�	��ɱ"���OetR���IH �h� �"J����/���om����h�e<Mя,=�RJJ9;�{2T~pRw�x�bھ��k�EgK���Ƨ"����ؽ�3N� (W�d�a�.:��� �c�ǹԼ�V�F�^�&g��-��k.��ŭ���\S'eP��6��3�j�9�(��@k=��@a��<���+̅~ضe��P�[���Mc��ˉ{4fL!p�Ь���X�@^�����B�n��q��SK�����DM_���@0$��G���N�:�p��MzH�DfP�#� x&���~���;[Ϩ4��p 'Y�PE*2�N@ނLv�#o���!n�c�V6��m`:�S�6�����
}S)�<=5�V�A5�@]���55�zr�Q��R߉q���z�E��u�u���
��۪���L�?A�X���[�H��G��wl��+f�ϲ��o�=�+���7�������ez�d<�HP�����b��_��>�^P'X,�$�]NJ��K�V�.
�s���n�Y�mŻ�tf�X����#f1��[��f�J͉!�ɽ��ȶΓ��m��dLP\_���7*����N�2ox�5��);ir�Kq�.��T��{Y6���xu�9MXj:��Y��d�����OGu�Vd�`wu*<���Dš��?̲%{N6��Ȏ��O�\�1BB�,��ʊ��TD ���L���?�ދ$������܏�p	����
K�!�����������
9�g'��aX��lq�5fb�����,�;L�/5E&{x�I�{SY����4l`\���u���cb�|�1���{�N����h�g�uma����/�wDg��r�>oQ�ѱs�U�-��m�@R��v�W��{fSއ��4�Vx��Y�B&뫗�gV.��
Q 5 ��J��׻Ϧ�}��?��g{0b�N��oژ��SG[(�E�K��K�J�B5�~�|�'�=;�ⲯ�D��U�#�+OM֥�(e� ��}񝳲j��"�i�;�]�hʅ>������ܻ�2�*��*�$&x��-؏���+ֈ4"��6Ď皠d�5����z 巟�S��Y�����Y�7FR��M0&��b?z���6�OuU�rit����2��'Zı^�L98{r���!��\x[���9|�@�wދ���Tz�Y�m\'���;R�nZ��{C���ƻ�0�`8ͳ�&�g�;5ǇaN�����_�׷��^V���P>(���A b$u	Ɨ)�X ��AF���&�fFG��Rb�Fy��O�
��g�ѝ�*��L���˲�6w6���p�K2G'�'��J�1S���Q�H�M_�y�^���襷�|~���s����CD��V�|�0��|h<
�_E*�S��9o��Cۀ5�����y��jk��AL\���'�a�����?y�[���&��O�S�UW2���_&(�jC~eS�M.2#ٖd�����n,�7�8�==�]>�$�O�I�Cw�i"u�����_�*$�aWH-w;L[� s�%��ю�ݰW�OCūf�E��{��eܸ�go�5Oan���T+y=w��7�m`��=�s	�>��j2��uy�;V����'�Y�O��PQv��#���e0�,	KN`�i�c���"Q�u�[�,k��q0kHXBb�<�Qe�X	)��dwm��n�s������M����J�'���0�}i��Gs0����a�cZ�Vh�/������C+��v@|�Ϣu䥔9cFz�;=�y�afg�"�۵F^����p�LP*�E2S}$�ş�S�R���3г6q����l�'�;�℩{��0�z�3zg_�<UG#���,�������>�U���?A�?��9i9�c}�7�� e6����p��	V���o���<;̸�Z�*fOi/��q,q]=��f��8o��:o����*1�d|�;�m9��_\�L�ܬ ���٩3�����{���@����
����WNkOS�z^Q��:
��6]fN*����n��W����ʖE0EvG���>��%���`�/�5��8H�U�KF/��;y�1[�X-�%ˬ�?�t#���|������	&��Z
`]{!����,"R�}k,��c�����ҧϹ�أn@��-�~b㷵���}�=ҩ���jl]��>�ٝ)s��w�s,_���D�����Bjii��7���m���Q��V���}R� U���P+�)b��(���yc���?�,���a��4�BU���,���OK�ݣO2��%��c-�BbNO��C�6K%��M�p�/���s9��+Ҧ(`�.r��e&�YZ�䕲�9�$VP+�aRM7����v>�v���}�.�:K�s��X)�8��Xp�7c�eխVş���SlH�������͸;;0�gh��k#�"Z=c#��'�T�ƽE2ǺF	M���4�W$C��Z�~��@4'9�k�Ė6��Q���o��]ђ�[u�2�.���B/�U��!B�{�J�-��S�K�a�zAg9�r�>)���<����WZo�j��
���+�CiL��-�O�@hҞn#����8�}y�1-E��a3���s�p��j&ev{%��x���S�}.nna׮�� ����b�4Ê�p�W��\���H�`%��Ȃ_������.}e�B�H�V�m#����e�z�4k��ީ&��|b�w�̅G܉��Q���u,�gcr9l<�4�+����5UZ���V���Ħ:�X�M7�'ceY��]:^\~�1���߷�z�Vƻ�E�[{5��̞��e��1OQz��xC �j	a��b�~�l�"�Md���8i��HH|ڸC�\Q �W�o��'\a@ ��W��n.}&�k�7�?p�T����u�m6.$ϯ` |.
壣�!\��D�2�hDғ�h׻l�L��[ϧ{�x��_n�&��zt�VU�y;|a��xl����̉�z�@@2{�8����Tn��|4�H�ۂkʀ��Ev:(!�m�!�'b��.ȓ�>4mФ!n&���h 
z-9�b1�RinZq�����ͧ6՟�/�;Xf9�Sw+Xi�Z-��Щ'�Zq��<rN>��m�!�O��hm�.v/�.�Bɤ�@H\�N�^��D8X�˕��#Mnc����T�WuL�^p� }�<��\����F�{7!}��W�yw�^��Y������S>��R1S����(Z�n�]�{Q�C��F1J}O8oA��M��Z�qB���o�<��G�CgbG������������;C���?B��I>��n�_�A�u%�r�T��ߵ�g��^�Z���%
b A�}2n�3my��*Z�&Zz��}�t��I�~xH�~݉>ˉ[$E�A�D!1�ɦc�T���x�-��jv6��ҾRA��\P܅vDa�ji�� ˜�lߏ��J�~��\%���{��㳦hi_�Y�<���q}�0����4���E݅Y ����g��Hu��L�R�ص��@޶�:�����q@�ܾPݗ�+�XS�H���'w?O�>&{���»Mȅ�����̅Z�V46�4{��oxۢ��,v9��zg�H��x�㝲����dֹyx��x�Z�=��s�(T;gk���{
�#���k3k�-u1nS���<\�}�J&8�w���,1P�.Z��kc����͓�:���A����<V��gk]tq�Yim��n@�>���e��!�Z"���7�% �����@*>������x�~ֶ��Gߍ�}��,o�8���F�[E�ە��[\f[;>��j=����;��#{Q�YY��S�W�P��Ivg����dQ��*���IN�_b��@;rR����f�)����!�,m��乲�g.��ҽ<���q3Y��D�ũ��, �p�3p�&�o�fo<fxoc�9�@k��\����AыK�1;�����ȧ��s���sJ�>��-z�����o1�W�)�%�k"�<�,X���Ք3��]K��tj��hi�ku��]�as.������èAˁ7���;Y*�s��:˦(euU��K�v�`�d�A�_1��@Ւ��?�~��=��0���`F�TnH��k���Ն$ c��GЃ�!`�48���)�9�U�`&7�W6��?c	8�>������	����,��UFA�عVw?�g�ȷ��/�D;j�dJߠ�f,+E���q]�����+��?���8A �)��zs�R�31�\ϙDw@�Ŷi���!�4UkG^���1�fU^i�t����/D�=L���r�s��_�	��V �p���	��0d7���D�^T�|�����"���KSl��z|�2����a�"`w��\�=��آ~�� �3g}�&f$^�ҷ�S���ImhY����wRB��8���&�&���|�������l�� H'�u�� ���Eؾ����l�k��i�N��ưND�s~��;�M����$�F�3wt��V=v����r��B6+�3�D�|�fY�=�<�z�tq��7PP֌7���X�^5��:^R313�K�y<QiOE���������/�,z��άi�\�@�Tqy�`�֞T*7�%";�]
M>�;�6t �|��5 ���S��{���6y�`/u7�����SK,;��뾒ܤ7/+(��{��?�Dҡ|��:/��J�B�:�,�
)��}�A��ol�F�d�T�����͠�K[�n+���qU���!�� B�mv�|iƶev���g������=���SFCd]�<	1OfPh����B��j�/o���¤ʭ�$�$k&UIb����m|Hl+ϟ�:2ŀ�]<1�-++�����Vw$�N��&��	�{����e�����2Jd~l�&��5�8�ym��]V��G�j:��\e5�? ;�+�U�3+��76��-�
�鳷��>3�|H�3 ��@ά���e�� �u���.�g��}�@	ܹ�E���c��Jn�j?�&W�I��uG9�|N^�d��:�'�-�s����3K��^����:i�찑n'�R���]�ugt|\2�fصT%	i�O��7����9s���a����� ��X=~?U�>�UIv{Hl|ؐ�Ns�$����D+��Qu49��_YH#d� �̙~��JEw]�-�\��3�w���^f�^�Q��5�YU�.71���;tSjH�� 4Jf(;���ao�pf�O�oK� �Z�Y���ѻYm����u�}�j��L��JJ�k1h�P�3�yy8�Ʊ^WK.�*�(wT�.4�x�N���XU����o��/#G��-a7�I�H>�����u�g�$1�䈴��#K;+>(5�x���&^�4�'��=�7 ]P~<y�X́1�$��C�O������i��mvCo�Rv�\ǒ}�X>�r�}�,��K�C��� G��	�4oI¾VW#i�h�;i�/6$^EG�Ayl̆z�4�{vf#CCt�;ב=e���t��,���&�ט���wȫ��&��;��죨��J ��F�9�%ݹ��][�p��R���>a����Ő��x�
 �"+@�7���?��_cl;�A�����J �((��z�vB�J�,.ug�'V�a�/h���/��_I�ț�Tr�Rh\]�0f~��ѝ[+`����Z�<l�uҔ��o���H"{ќP��%& S:�&��� i��ʲ/ҫ�+NGK���m��7�?���ǫ�Pͣ��|���>��{�,��'����I#���k��`�BsH.��0jHjϯs�[���Dɤ ���b��p�)���������p�]��(y�dj^���8^S풻�Ms�����G3�|���;J�8�vߍ�7�h�*���)�z����r �a�[����Ѯ%w�c~�E[�ץ.�M�0�)CRi��>	���^+��}���v��|��F��ZO���Rء�3`x�;0��ul͞�U�o�~��	���ů;��4���\KƔ"N�2r_��>�0����H��TC�o��'2b�*X��� �`O�^�,� ����;
��گ�{䥺��n\���X�^I�`A���Q�(�,�f)b�p�����H�ƌ�^�g�[\���uu3&⬕ŝ��7��~���z��g>2\��q29G4���g�6���2����2�+$J��KX�'Þ�[��m��7�
���������;�a�7U����g
�9-`2���˺F�}����	ӯ�VslqH�g�7�q�ˊ�+,<�y��4T=�J��^�E�O��$���]T�M&�O�*g��N��<�ip��L���d��[خ� �7]w-����e�ό�ʙ?���楨#����S�G����!��ÂU�!Rz]������� wDD<��y=R"�d�3��c�^'��՞B��)�S��F���ڥK��Mb�^�ǜ"�)��c=|{�ϕ��.����K_���0�ߑ���]���b��_��W��t�6�шꉭ�5RP���tuER!	�9�ۖJ`0 ��e&�*w$�&U�����"��J�"! }���겡88�-~DR�A�#���C�|�D�����q�/X&sdw��s�7h ��8�+�O�ł^��6ď{	L v(�3�6p{�P�6ƧEVZ������T|A����b�>�x�S$50��)�6^��e9��/����k�J��S�Cy�E���0��𤆣A�|8�m��M=��X#(ѹ&����хd�������خ�&m������E�>'7(�y+�SR���8�\n(6A I����SO��~�ų+�����G�!jo�@ n� �u��('{`d�V
����e�uv3�y�O�N����b��u�/a�Ⱥ��	(�*-�L*KKz� ��x� �H��8�.�=��HjKj�(5�Mq���a�\QϨ������Oܶ�Yu�f�$�L���R����M�/�	[/;_-�N)^uqѐ��d�w�T�Ł��];ȭ������y�_��ǖVV\��kt٘{Z��H���"_�M�y�އߨM(�"��y���?ڌiVt<voLpYWCq(}�w�۸��8y(���A��32�h)w���aЫD�Õ�V1rYr��*�r�B��P�g�]�7�!O:�X� �h@e~�G�`���o
��L�vrK�����e��y���H9a��Y�_�C�0�VE�^�����΂�W �W1�i ��N��^�G�x[5�
�ܐ֘D=6H���`s����$D���o �$����
���\�S��� �$�r������6&�����a�㿣(E^(v���V@T�-�^BA�?��.��))|7+�(���A�~�k%|y ���s���s0Y.�[�w�ڭ�RDZ��$k�E�X�0e�;z�f f�Z�?�EtX��G
�!���̌ڣ_5r�۸�ءE���@?@��`�7�R,A1�8��W�,600\���f��?����I+n襵42����p�Y�L�~����U�3��$V8x��Τe=u-��P�M��Gփ`4s�+(n!��Wo�3j��D%���ݑ��g���{�zmY���Z>(���+3�e�9�-=dF&&'#|t�A�u:1���}������!Ԕ������$/�6�*<4}bO4�6સUI���*K���VB�^b>ڸ�:�9;H�|\\A��h{�I� �0a�r���J�qDX�f���1� 8���mK# \������	ʕe�1��k�Qd���-��)
O����?���:�`���y��1}��E,�>���8}.(��_)����y��~9���h�krٓ C��?���n@��a��`���W33=�w��dǊ�k��4��P�o4�kտ^��a���	�-�=�a�j2Dخ�zW;�#g�O+��n��
����N#��������0�`�ѹf�T������B]�)$!Qgt~�H�?�5U�S�x�[�>�_�7۳��y���1�ѹ���4�����Ʌ�z1�W;"^�����^��'���$�M�����ݡ��}0�f	��־���%�q�p��nM����5����í^��GW�L;h����Lv�Ѓ��u��R���R>Q��V2�o�|m@/l��;�cԨ_|�`����m��o/�}���(Op;|ed�gKpAP��H�|�{H}�0�;�7����J��Ҭ�����G�?���bR���ARK��6�7��A`�A�5��彚����!�@$�O�]�4_QTX���h���6V7�~K��zM��l5a1�3�]��U��()/oJ�ޱ�`3]���k3>����֙�h|�A���ϲE�ܟv�YuB}�&$$v��#��K����P�]���$P���|�ڈtdO*{���??IP���N��ۧ����Լ��$S�Q�N^r�h�!�!�#[�V���ʫ�S�����w&,��ːG��x�sIm�\f�׼E�l��Ɯ��ęO�I:�E��y��-��ӺZX������oM��F�m�c��_�,h.ӇE�q=e����T�0�W��(F���WW-n��sz���,��:��C��x���
PH��P�+�T������+�7�����O��K���7u���,O�d��_|���-�Ӂ@�9��A��RnB.�g̿�XK���&!����2�1EOEr�X���&�D�zn�zoc�.&&�ؼO���z�=w��̆
�i��ih��ޙ�ʐ��4R?ٴX9(/��T�a}�ɷ֜%��h�Y��Uy�p>��ߏ9�!�����]�fb�:?M�]�W����xj��(>���40d 1ک��)J4����,7����Z�CX�6�Cq�C|�AF��%���������ah�L"O]�idHa�v��V}}�~[Z��hBt_U/ꁡ��N�)')nK��1�O[G'F&Q�b����9�(�j:~�I����(�܋�ݲ�浗�I�E �)�(�x�&���iZ�s١���f��Ml,��5��,&��4t�;�p�O�/��ls����O{�0�����f���9���:��A�Bs���(|��/I^t���U�[�W�镣"�)�z9)g��>Z���4��x*%�2�@d�*/ɬM�\NN;t�Hw��)��L�1�� ��iu���|z�Yȷн�
�\���E�"IwF�Y��AH�\?5�A�rpD6�7�M�w;�!�򾖢8��:��O/���H7sV��o��:p^�g>��Q�aa�� x��u�B\��� ��ѿ��w��q�K*ɺ󺥑��2���oi�A���+� !�!�p����A�S�B���[��\�I��	�~OM��8�Sx�6���xc�'H��V8��],���g��(l�;;)tDFΈ^���]�c�������mE�_}�=
ՠ�>���1�d�Q���P[3���h��߹ŠJ� v���y�;pժ���,Qn�2�wٞ�(_��l�S/w�8ϭQw��M�&��`q%�����,�����(怶�0�w�W�C�O�5y.vŝ�ɲsD�PE�p�������g�������a�d_��QWQI�%�8[�l�S᯦����'`h��{@���Z����O���7\@�\�A�I$볘�-^(��
#
׷U}.?[ApY-٥#w�<[�7��A���Y�>�Y�_X(!�d�꣘X��X��x������^E)�5��4xN1��0_N�T_�|b���긠6�c�u����O�%�z���n7ڨ7�z�
�E66ɖգ���Z������8�n���a�l���1\���s�u�E��%��@�?���x#v?G�}(x�"Ȓý֕U$���HWnOL���	��UV��1���6���;����v�}�cK��3k���!��j�1W�h=~9l������" ���FK����� ���Qi	:��[�9�%�����X2&���d�3�1~u-�#���Z��@H�=�u��[�Z3GH'�EM�ګS?BX1�������2Ł�������~��}V��PI>ǰ
֔�'�����'���J�[�.��xc��QF���0U�i��U�=��-'�y��k�z��\�߈DrR����w���o-�[�ֈ4]JbkD7��	`�+-P�s�'>�gdI�4k�&�yc��a<���q�_"^�S��Y���Q�{QA�1 ί����Ț�ONUB��@��Q w[�>��6 �I>�M�|�b*���Y��O�v"�2��;`\tTӿ'�f[ke�|��?�x�!\�5��cӋq`��: �;�Rf���s�����	��m�}ŉ�]���M��v0";�d�-+㬝�EqД�P�.B�)F�ã~�qWid$ѵ�������]7Ko)�.����G� )8�)�ܮ�Vey��Z��&l��}�����A xa���_����#�J��h�cT�+v���T��:g�U�άm�u4� MzLE�>�o7dS=��v���ҹn�Q��`�!��؟��N3��^?/y�s2>����?�f���o{������"+���`GWCH/Fj�����r���N�vwι�Q��۟����
��z���������m�L׿Rx[VV��a7���<���0������F$�����&FF���GDY�ܛ�`�Iq�'�z�r�ļ,�� @�j��zL\��,�����f�Bc���/.j����ð b��e	S-9�tP����K�����m9�Hgff��lk��ʶ���3V�^�w�ns����I6���bAE�Ǯ��ζq�%E(Fj�x�{��13xBohB�2�mXY�;
.,�ib�.M��'GCI<ZW�A�O��<|������n6,���:�:�ʵ[�}��y�c���Ob���e��z��w���N�E���.ϧ�^��� ��%g41��ūH�L9���*�[K����M����Z��
����NF�r����п�|�6��E'@K}{��<A�iz��|ʼU�m�Z��	%V����7<��M�/�W.�{*"����;[��T�� ¹���7�E�����T��;$�v�䗡��	l�c��~�%Bz�nb!��i���w?�5MQ<~���*�̎rV��N�2o��#��f�T�妦�jͽ�Bf,^�d-�OO�P{/��k��15l%�3^p����4$�mɍlx'��÷�.�O�I��8��5olll`�?��:o@(w�D��oͯ�|�����7��f��1X��;��CV���)x
[	9�[�nb�_�U��#V��E�d��0'9��q�"�`u���s�b/7���<*�b��S��O0]u�E��o�?�hͨ�)>�n[=�p����7��k�B�� �,�<p���Wc�it�+V�̍R���S+���F�{JDb�wu��V'��ӓ��@���$W��c���D�̞�ӉJ�`�ҩ!b� ׭�m�G�����擗��#V������f�Z։=:�&��W��i�xV�3��H,f?+�d6$|�N֊���D���FR>U��|Jh���͜�\���p%���K���A�p����6h��n�>��Vw���=��r{�����Yktp0��>R7�IV��Ӛr&��{A�Heig�ł�&՟xu4T��.�?��L�T褐�!����v-�n���u�����k�,dU�4�L�(MΏ��Ԩ�QgR��Ǖ_B���0�$�l�P���
(C�e ٝy�2�\��ŏR<����I���S�QW	�8'�d(�hi��&l�~KF������1�Sg��n��7���t�RϤf{��B�P�f�ٶ����i#K\W�9�_epы��^�a?N�cxݽBWY�Ǧ�$� ��/7Ja��6�5��&�)%T�*A������rA�$�]�S=�'�OT����Ky7/�	V9 ���# P�����[���Tg4��� ���!b
n�l근��'6�jԵ��/�dE�,B�U�:�d�*��!^�V6w]RK��3�!��g<�����;y�'�g.���}�o��3tO�qW�Wd0��xLWr`��m[�:����A����������p�;L��x��]zRQ�|���p�������TFyyy$5�Z�I�`bP�}8˨
���9��9�nH0���j��F.P�b�S��`Ӈ�d?X_�m���c�cL�q�6�7���ؐ�ɓ!������ٕ:]q�����R���<Z��'�l<Z�f���+3#K?�����Hy�tR>�L��m�#�^�7Q>��s�D��O��|Jl,�-ڎ5l&��y����˥��(Ѝ�*�2�M�VU��%���9M~P��brf�ᚭ�o��uM���$�J-�\��/��I%��;����F��_�gZO��s�&���Zi�.�߸�j)��9���&$X�C���D�5U�=P���9�/
"3 �F^�8��J��ۚii�=�v��8k8��E�)�/y]���[���T��	�j����jn�|�2��-��A���p'7ȿ��o��"��̞���0i����I�x]�`;�m�tv�f���Q���_g�`33�H�����dc�䴆��Љ]
��ߜ�Bjq^Gb(��Ǧ��EO�B�)��T�J�f�t�h��¿^^P���ڑ
��O�!3�ҿJ���n][D��ms}�H���-m �|��|��n������E�<ɯ��^<n��@�{��$p7��vA�y9���o	�f:�\ܞ6�?	��2ґc��Ԓ� -Z��͔Rl~p۵7�>�?=��aU��߹�&.�hE)u�ܻR��w��L�?��rݘs��0��*X
`!������DŔ�MvA�%](�A�pf:����%��[R��P��ޗƿ�������a�i#�&1.�D��a?Ǉ�=�Á|�N߬�?�zO,n���o��`>V���Kj���c��|��R���Ѝ,#�7O�cs�u�ew
�N�wTthlaT"��ed�8�vf4q�rb'�9������X8���"��z	������i�_[����J�����N�*	���b��X����S�����H�=���!��O�8�fp�PM�D$u�[|�K8W@����v�1<|�V�j�� +�Nb�o��z�''��υ��&@��暛�/p�y�wc��9�ѳ^�Z�u�o;����<٘j����mD�Re���[�Í�������/��?m=�^A\?ms�k+��v��ޣM����g�n�6j'�n��`�=�;�~E��]��탩�|p4��@";Vw�,Z��0��4��Fn]��W��n�����.\"��A��<P��4_&�괳h?iY^��W��vF���/=�l��s?��56���A"��#�`w+��ls��v.,�b���T).��᯸^��y��c\�U�F�pn��bag�-�=�	�۪Wz�JAM��'�4�yuu�>Z��������,�_M�����K�@?Q=&�Y.]�n.�Zb݀|��&�9�7��Ul(��(�~A�#*ut�}��/v�!g�v��|���%�q8�=���ՠ>��`l|��x�o[`��M�߇⁖#%L��H�|3��<G!����W�jxS�r���N��Z��3Y������c=?=��ܺ��������"�X3s����|
�q��+M�Q!��aA�MI��^����,7���էv(�:oѧ�7��?��*����F��Fi�����A@R�n����F:�[���k������_�,]:.���w^�����6^��q���-�ȓ�L���x[�O��rz˸��2�d?2���7~{�4a����?�΍�vM�{s:���,��638663Cy�.S��d��1�mQ]�޲��<U���T�4�A�q��7A��p ����D N�v+>�.��[9R���;d�(�cV<�Y��<�#iM��"/y�O
 K����J]O�`L��\��.���%��|"����~�]K��o;���OB( �R?�
Y&��'$G��H^��u�O񠓕=����I�Cw8a>�H^�_Wr���`��O���������!��=�L�l���1��W0}�d_ )�oH�(ts��ևN�1 Tm��M������~�T�Ԙcj3O�s�������麛銤P�m�i�d��o3i]D�\0����H��z�����_!$��f�1&�.�Mw�C��i��nA���ڑ�_�Z�S|6 ���XGh��&�ԪmA����t�9�s��rP�75�8�R��񈗧���z2�5�m6<��Eظ��j�A*b�=,�Y����UN���@�iX���n��q�U9���mG�o�6IEfϥ���8���8��d5n�Mk�du8�7�v�(���ܵo�%5���i��=#+��_�q����jh��7JOő�Acb�d�*s/�|X<�p�/��n��W�۝�?]��+~��z��~v�s��җ��~�S8c���A�zu�r�l�|xHT�
�f��d@����F�V��}�>��ϸ�_�-���K>B���iE@(�,��a���9�XN�����$F�&WT �ɻ�$)�j9nT*,fx���t�sz�m�i���B~w�����M$Q��%'I��v�E+�f(7��	K��N.���jW��_Mò���sM��n�C��l#� YW ڤ���W�ހ.���ܵ��&gF6�À/W����Q����bc��꙾�ك0��f?����� �j�^$�>�W<��,�s&���Ej3g�/$v��z�}$�y�Ű�H#ޅ'G�$�.�����[eX@�ߘ�۲�̘�+��;�I6�70t�����(� ��m ,6k���
�Tၹ�~!�|(���� �T
o��v�������j�-w��OQq?���g����%�W]Ŏ�p*W-���'�E }��K��#�F|H����z�q������)p}��to�����Q�VqC<o��"�=P�P�O*��C�,�|�t�c���\!\��@���k��p�q���q�1OM���w���o��b3�K�O�����5
�xpB�&8)V���nD�(��*�?f9ܹk�˜MJ���yJ��~M\S3i���njn��w^9?�>��E�L�-%��a'{@󇮬1�9���d�JR��j���+d�`zjΈfJp�f��Dnq�45"�=͎k�=�)�Mڼ�7��/V{���ϕ�6�ߜG(��>�-�g#�宍��������ЇP�ܮZ~Pz#t��OY����Aj�W�����wcG!P���X��ߺj4����-�g: OHݷ�&�>��/Lwy4�X�x�dZ��\��0�͙��R�b��x|?	�q�q�����=9b�<�ܑ�o��fR�W@W��xivQN1�h0�����N��.���	]\���>L�rr��|����Y�w�V��Qqt=T��\����'�N�""(O"��G�`Z ��%_������('T1�@5Gb�Ou��`�Χ������z�"_6���*H�O�����WH��#�����T �z�<'��Th0�OwqD����jt?3�z��V��ErC�+�s�:A�RBZe� ,u��F���4��ٓ�}�����(q����yKѻ���W�����/d/�4I�0H?1}~��}2}U��+Ǩ����t�K��RV ����4#�nK���#V.a������:4I�bv�2&��ݑ��;��Q~����u#���]l,,��6�$yDT�XX����L�]�Kqj�ވ�8��W�|���b=�ծ�9��JK!�h��RR�V�ϒ����G�
C&�o�3��j�y՞���@?@�h.�%�"h-����f���� y��n�K)G�_G��?��0�x�x�w�y�������aB���Kc94ߜ��T���ᆰ�c��k/�����;1��'�]=[K����M��F|�j7�58���2Č7|��sF��^��K��1�Y�-J�w��E|�n2XS�n7KV\l?!��=_�F���F���ʟ��j���2���I�L\�a�����'05�0N��˛�]���f���¢߼�������<���NQ �R*�ǭl�Lι_r���;}Y^��}U�i��q,2������%d`,E���:�m�(�{]0-�1��G��a�'E{�TC�4K���fۘ���Y���࠾E�g��#�-���ŕ޺��s����� ������Jҙ5[��)/���߯<�k;U�.%L�<�}��L��o��0���#����
_懩X$Q+�Μ��&�����F,q�1��(���6�o���YSyyYֿW���y<�F1���*�eZ?1��pgo�$ ��g��G�o�Q����籂����j�V�?v�Ȱ���
����M�}�R�������ßIs+�N>��?��4e�0G���}��C�F��qLDI�O����&1�sF��I�?��~
O�)�wL�+�y���Q�2���Y�phZX9>��Jg}�|�`���P���7p߃��νؑ���R��V5��屑�J>?�����X揟Q��$ỻ%�}��O�h��6��|On"�����x��(aE�*�2�	َ4	�<�XcY{����x�{A����t�e�N=j��Ň���IL�ͣI|�*sz�\펡C�s"zq�ý��|%�|y��~^���}ɟ9ř���_SRR˖5���m��TR�3��IK��ҵ�k�ѧ�����.�x��`��ƾQ^w�{AF��]�y0�*�F��~1h��j���dQ���>�������C{Y漏��v����f�(���2zS�2����:��'=M�M��t��3�/l��X��q��r��\ �_�D)bAg���=�q�@xCs�#a�{�v���_AA�b�Hq,���m����E�^r�-������D��y� �_)�k?��u��s�%�=d�픜6;����>���o��{�<.g��>*�mcJ��.���w~�ttI��5#^����sn���Fؠ@�IN����yE��&v?�k����tէ���C�=h���f�S���<����0��4i"���,�R��e�Y�}{�&�� �9�J�f[s���灯HF���O�kr߯� ���K~;u�P�R���^G�`A�l-~(��22�%i؄0�\�f�K^\|����-�34X�2N:S��GA����V�ߗ���ْ��jV�u����Ӕ��,4��ru��E��=o4��_Փm,p�]��{,�z>L��p�)3
BFJ�S�m�9P��)��Qq����2�T�o/�{u��ܒW�� Hz�B`�vh���M�Q����SYָ�h$M�_8��(?Mq�l�����}_�jFz<��?3�њ奚�j�ʒ7t�rR��I�Q999��"D?L�&Ml�W�IZO~�X�w̮�Tj����� JD���\䫕8�:͋mw#)r5��I�i��d,�����?Xiƽ��i3���m��|G8�e�M��������+�aE�PA!H(���ko��ޞ-�l�ޮ�~�R���sr�4�;�Y�wo����|v*�l~��PT|�&Ud nDig�q�{�1�
�R�h��6�	�`�R�z��6����r��ܥ1�Fln�
�	��ң,A��%c�$=�$�ޏ��B�<Nsㄒ��L�;4uמm{�Q�hF�)����h��$�)�d�;��q�!�j����~TJ�0@A��
O�|�v��c��V�=�Y�0b\k�1��*ϥ5B�h���-.8�;n�x�z����Ѩ��m�e�{�<��	/�񌇚��$��W��6�֋��fgW$9�ֳx?��2��Y_�*�rb�r0���.�ϾE�<Ŀ1�O1j �]�O[���U��ip^�֞����F7}���H
�](	p��H�$S�K���v�����U�2�ù��0V��T�i�"�UK�.VK�tkL��O��j�j0_�WV�I��w��I(w�,��1
�*��EICw�y�Y��]'�R����!Up9��ay�5�[�a�/OG�ֲ�`R.A/w7�UU�.6�!/���>eǔ�F��Y)���k��������-�0I*�^�vJ̆H	��`���I� ��w`��F�y.�������UʀQ�9R�{D�j�ڄ�^c2�B�\[�e�����-���UK^��
�E�q,�$���r�����Wb0�Z��'�[����i�����6�� 	��PR߶��	/�FK�����M)�vq�[����پ�������zŖ��r�a����1���o��#A ����Y_����Th��
�s~�!$D��/ ɂ�}C`tA͹�Z�<dr }ȧ�e?fJ���R�X�V�L{�o��-���.AU���:JV�<p\�+���F��Zr0:nvO����u����Ɩ#y��C�H�XoGe0��D�Pb�f~�ϳ�:�W�ٱ���,((�N�` Mg3��7�s�d�2b�<��P�	��IiD9 :��o��x���d��9qϳq�n���u3��D�ݤ�R���M����!ҝ�.$(q��W(i�[  D���*���^��0����� �X'&�C�4�d��.�*���`ij�u��֙���̊�����,O�����m��A�)����?���.�|�����ԋ�f�Z�(������A\��2��GKY䎚Z���Q4��0@�f
T��Q�
n߮����@\!e�����n1�s���H�����s'��h�1�Y��@����I��ǂ!��%�r�BD����j�]k��6��J�殘`-�n�J��N;�ݍ�n��&{i�M54�>[H�U2����f����3)a�?B����<�w%,�p��y2ֽT���>h���Թz�L��Nl�������{����T4�5tjji��-d��죳�|���A�gV���\(�1F�*Uk �� � ;���\�EmL�?uc�Z�C�������8@9���[��nK�k��Ic&�މ��@w�'db�F<�=m���r+$��-�hA/xD>�ŉf;m�2Dܮ�����v��>�i|ֲ��[�^�~;�l����H�y(�/���%�c��E�S������ejkP0�`�(P>�K������ɶ}NJ�xϚ����;��m0i�F��A��i�|�_���Lq�P L# �o�����o����إ�43ϯ��x^e��4�]4c*��Z�^�ڧ*;y��N�8c5�kq�v��~W=�0%�bT��v�����j�"�����	X������gy��uNB�W�a�7^�++3Q��.���%�[��傐j�t��������v�fLhi���#&�����`�%.M�:�.@�E�	����,�����k���*3�%]&�^ց^���#p�\�L
s��T����9���4�F���� מ���`�X8���m*38�q�e�#�CA�SF���r|q	�^%�MC�K ��N�zbaYFǋ��`�?",�RDk��E��`I�y�]��/{��$�������E㋦�C�@.N@o��/�th_�2��&-��k��]��
.;S��tU�h=a���F�@/ť�Iǖ��E" �&}�)��C ���j�M--cI|��w��P�(����N�ͧ9&��B`L^���nQFa=�|k����[��»@NL��u�l'���~WʓX�$�1�{W�ly�(��Ic
����@A�N��}9�`��?�oK������u��*�Woٰ��|��L�sk�]�*�Ἆ��ԩ���s*S	~�_���m)�w���U0�z�@��OcD�Y�Q�r�Bvm���ּ�f�{E��w�������L�Li��`��u�SJ4�����/�	JƝ�wG MP]V&,*����̪�XW퓌��Lᣬ}3�V^���ӻ�ךo����Rڴͬª�d�L֠������d~�>1v( ���XL��`>*{��n��j���{]ۻ�0�q��9�L�ǖJ�#9����~�q�Mw�L�����.#�W�%��͑�@=88X�u����Z�w��k�@h]��;����a��5�ΦZQ�]�#&Fm�y������,�������eDt�
��ʲ����	諁Z􇬥ٽ.��s�WɋL?I��2m7~��8��y�R�;�}���+���&4F�,�rJ?R�Ѭ�ш���c����bR?�r˹��9��6$d���4�w��O%+�6ݤS\��"P�Y!P����U��Sv7G�d��g%[eU�d[����+���o1;U�5q�����l�0�8������@����f����sٙ��5ũ�Ͳ� ���c�˳���9X&՚`Tm9�d��iĻV�͕j�r�=j��	$?�lREFo�eR�o��O�:�xq��b3�[[����'!��=+]�{�ݛ0/W8�'n� r .�M���9N5nRR�Pu�aV��=t�_:����&j6��#M�į��
�!�WM+c���3Y4��ՆT÷Wq�|s�#���PN�;��}<�Q�es~��7f�$��+�kÛ���h�R��f�~(E�(�˔�ZllY��F�'��>F�{ìc��z5G�?��ٞ"���_�v37�7��6������칰���c�^Z�(��6P(��x����=�R'>��(�ѷ�Mթ��\���2�B%��-����^9��-c�(t��z���˳r"W.�=M���5��
����ˤ�'WW�jL���ݦY���Z�AǕв^�𘲓�3_���������,q�u����������W�C�S��
�ȗ5m)���>�Q�������)1��11ہ�phf�QZ^x�9U���5P�o�i��=�'���1Q"G���Q\���FP�:L��~�3�����C���WyI��P�
é��?Ɍd����[X�����ٲ�U-���� �u�Ar�X8��אC�§3AՖ�v��E�ZI� Y蝇��da��Hx�j�ߓ�FG�BX�X$�3����J̆�<�Z�tI'����A߬�O�*y>��y��L���������EZ���N*��!�o���s+:����kH?`S=3s�Ͻ�jjYEE��XQ.vJ&�n!���36B��.ξ�x�>EJT��;濧�U?���$����k�[���F[���F��p��#�L�~�3�L+]��[ى�);�Ff�}��%�(%�6f�*{*���)��v�U��i(Ok��=�=I''�8�d*�\ �u�}n^��`NI_R�匟~�Y�-����>[.x�;H:Y�~��[�y�V�z���Ū{i;06��F��W��s���X n���w����U��&d���'TSS���c��/�-U�F��T����l��A�&�T���q�WRӊ�d�+��X�o���L����Ϩ��[��
HY���9��9�(1��z"�kᗬU�(�슙t[��~�	�-�R����y��[ -��D��5ߏ�b���i�r��>I�Z��f�j/�})� P�bj��S��5���B�V�a��ϵ]p�����bl�w6&$��}��E�[��#x\m����CV&������.g_��">��2�jW!ny�T��x���H���m��_��ſޢ���돦��`������#��'��A�jʝ��A5z�.�{KZ�I,�_<���ho��"*�5ٷ�ɬ�<ܐf��*T��L��[���5ٸ&�)fՄ������+�b�||��������Qܙ�B���`� T�"�h(��_y��+�դg���j]C�IVB�D�'%2�7�7Z�҉�ߵmr��ԊV���`��31��9���X鸯���J�o?�'*w!�\�}ꩩ�{5�;�x�~�����G��o��)
��@W�.�@��c��#>^����q��A�$��w14�H�[M��<�Кl�!�6�6}�;�sp6q�lR�0��;��D�6+J�k~�-+Zp-���Y
~|ߋ"����  d��,�>1���sqP����>��@Mb�b����F
0�g{�����ԅ�������W'�X�ړ���I�����!���if����'|��p��\���2����s���LB��3���*` CUՅ�$��<K�$ٯ�zjT!�#Ru��U��O�K��j�ٶן�Wp�Yv^wt;�ʓ!*������6�

\��r���k��0�Zi��)5Z`�/��������*NGA��Xs )����/݂��?�bs��t4m�B�d�{��%|�v�3J�(��Ѩ#�����A�qӜ��|���5��-��E��9v�`z�F�ѩ�����]���	����7��һm�C4��R��^x��HƱv��+����J��&K����>��J�BHWQ�E�їq�Z��j��D���b�cnM����1�$����6��$3%?�ƫB���h�����"�u�se���t���)����]$��X0���T���+j����5�&|T����.��(����"q��λJӑ��e��\-N������\֤c\��lKY�ǔ%}�o��Ԭt�Ӧ������'���_�W I8�s�ئ�^�9:]�8���ם��B��ȊP� �>�9����Q�ԟ B�d� �3�aA��q�"�|�ڭ��*�l!NĔ�1k���0�n[����c�"�OW��8&�2W���^:��V>��T�:�Ζ}3�`�GjTu�5uGY�mۦ��,�b���R�6R%%��妺T����B�|ǆos�������{�X���� ed��ݢ�U��17�<��m��y�����T��[����%*6�=���#���9���p�b8M��D�<�e����U{�Q��9�b/�7]��bȯ��-���^�G�W�zM�3	���[�� ��F�F$L�Ǖ�b����H�zj����������G�]nx�|kxg�r�]ʏ������gַX��$�z��ٚ���'���5No-�m�v�	N�m�{�W���^]�Р�v����̞��zVbw��Up�;kY�f]e*�IH�sNP����7�S<��eݑ����|s\�L�� ;����`,�	���X��۝��޾�2�B����dm�s�l�3�IU���� .�=��L��q�S��7�{�)������Q_�%hx_#f�̏Ǜ
�䳿���:�:t{e��Cm��<������xafE$�^7|�ձ[�p7}�8;��'����j���O�G�b��=9���vI^��d�4��8v��tW̷� <{��N�C�G )I y�����Și�������aI7�Pμm<�wOޮ_�â�Yo�ۚ8W��>]K"���:YWW��!����
�nd�����⸃�Ƴ��{�Z�J�m�T^�Oq�[G`�m<F�ĳ����]m�>�R

������hj9��	j՝(��߿����q��_L"�v7����Šva��u��mK�D-�Q܋�Ϩ];�����°���4jW�H�S�S�JaoV��:�I=��!��3^,�����z�Z����·���OR���U�>����6����a�=\p*V;����r>�a9���n��(����]�XJ��N���U�a���#�_@ r������P��%PqaYY0�����{˷2�\�..�����{��N�J����¢"%On�V0�ݯ6D���ܫ�/�����i��|k��$��G�����=0"J�oh�d��/qҽ*�Zj:t�#�WW�]�}VQ}+Y\�`��p�K�n�f�ƚtA&\)�,�����Gy��́�����s~��]�\����AQN���$���iE�����5Ƕ� O�M+�8l&��:}���g�V?�?�ZZ.9H�Q����Q�y> ���U���#�8>�Aw^��q�pͼeqB�4s�F�<�#@X���Ϯ����ib�b������%j��4mi�:�vO/Fs���o�F2D"�,f
�xw��� �(�{ƈj��V֕�T��<��_n>�Y�J���My�!S����
g!����h vs���T^��aLW����ƚ���^�[Xd�t�4� �2USr�w%#o�Z������sK=^���1s��>ā��&x�*�nd��s�	���F��%lv�ǆ�Hî�kJz{����bp�9��GE���I���(z���"��^: ##W�O�F�����ǧq|hs��@w˟�}�OX�
�M��3Wt��0���|�Y�<%jk}f����:����lq�N�c J����)b��
?_�/����x�FH�����]���+��J"ILD՘P����`q�+�J�8�5�x�5H�oۍ������L�a"OD�I"�b�#�D6���n����N�'�I@ϫ�J_��*����
D��hڊ�o!�x?9E�j�S�	9L�NUvdZ���_��B�S�����L��><�eV!CJ�j?YZ2.��B����$��(&��ݻ�_��egSN�����~�/M����cPˬ�?撧��	'B�gX1���% ��]ު�l�����(�\�a�["��Ύ����?o��\�����==}P��TT��ɸ2�fk��OzN�7��Ȣ�����>��M'q|���S�.ʐ���ŕ�.����� 01��//!�^��:��/��E��`�I���*2���V��jp:������g��$"*"[uZm���+�{���n\{��=I�s��6�&1l#ED�&�w�w?�}�߰6�t��'�D��O0 ���Db\����E«�?�Vd����&�1�n2�'�7��|*�-�C+b��tKD,��g�.�OTG��-�����ݮF�W�59�8|r66��\M�}}��?V)ޏg��������t���'L9��"I��X�cb���Kʁ�&�WUWG%$,�_����������.�t���D �(+��/=��h����2�&L�p����k�����+7Ǔ��� �����S���0H��NU`>=Yq*��x�r��#�����B�����n�ؐˡD6�j���łۅ��R��
ɺg�)���Zt"ccq/g1����""�gf���7.�'y]N�A��O�AA0?�1�𧮲�������ۚ���9��;�/l�]z�##�0��#�{/�"\�&'){�>]����������6E����`�d:�h��?ѵ�_o'����?�؞��B�,�>��G������6�]�ķ�&�Q��28���t�������!��ς�K(�Ś$�sr�(��=�e?��$1�=`����~��W����!�&��w��k<���%�2�@#ڙ�_���
�<���p�Xg8[�M�lܱL�b��I�K��1S�x��IK�6X�����&#���f�� BA��]
74t��Bl�[�u�����t��w)ij���vGҀK��ͻ�O�����Y��___wي�Ұ��@�y��N�ޙ?M�ō��[Pn�{	��Q��)�&a�l��b
0�Qh�0??���Ҋ�RNN\��(Gs����� ��b��!@DD�]%Ds[���M�	�	QNN�'�\Oq0��6�D�{��߫B�L�����s�ӛ�1���&r��L�G��R3Xi��A���p�b�����_�d�f�����μ�� j2�N�6O2o�62Z�FR�R�q���G݉��(��Y�է��N��X�^�&}�l�9���5��.�iθ�u"�cb{y�����~�o�$�:�t����x�Ֆc��AFDlϕ�9����C��[�.R�oh�濫H���cs_�,��63���l䉗>�;�Uϛ���!�T'l��FK.��!���c���-: hjkk?�p�
���ÔOb���TK��'��&���峏R|^��B��u���:�K����(UK����%�o�P����%������W�Bn��k,9N*@�����J�|G��p(�a��幡$~`?�)V���2���h�����|��3��Y�a]�*h�m������9�K�H�{���ޚ����T��R�[�v�u_iP��(�.4����H͍L̀��-�1�L��W�H���%�[��U6�8*Ѳ���6��6�ቅ�<�+o����"r�
���u0��%��$ִ�#*��~o~�S�㮢��V�.��Z3��>.�f>�T����Ԩ4�K�8��1���}�wJ��~�
�����"��U�r@Mg�Y{�:}m��1�D�^���V�~�aTho�weC�@0�2��8u��l�PL���@ʁX �{�.�˴�g�[������z�%���$��L�/�������$�RCC������-���t�$�e��D��ؓ���{��	���� �l͝8�T��G���QPR�'i��o^�J��:݂��-҆�To�'R~r9���$���ܙ��鹙KyT�À6���}~Śքc��Nnw���a|7ޯyЦԇn7�5��ڼK=E�r�^��t�N��Lm�
]�Oc*��4/Y���4�Ȳ"���·|=�d%�0�%�S|@��Y�p���n
�Y�����Ŷ�q�w�1�cmr����Dx�\_F�$f��I���&Ii�����uInN�vJP<��O/�7qGGGHY�#����84OP�}�u��f�W_�o\.�yΆyV3vb��J��ʾ�Ђ\j"t�{�]/ƚ�m"9�npT��45Z=��a"�8�*699i7�TWh�r������ֵh�v|��aK�:=FUU���:�{��&�oQ��?��.f��	flH��7��2v���gO����/�z�֑��=b�my���������&�\���SW�5H^�z����7mG��=��5*�Y�܏�}w��M�g���CA>"�xrL\�~���I9�b@�4J����8f�{)�]�c��,���O�ߌ_Ā��e����j����޲��j��Q�͵Ũ� ��q�)-K��Q�o2聓���emO��mH���#���M��
#��^G����X-3�h���O9�Z�Wf�ƭq~���eg2��#��l	��/���T��Q����WX�7��Po�����s�#&{8i#��VUt`i��O����'����ٞ�t�&i� ��o�������c��|~nϨ݈)tM��z?�v��&��g��ED{�ǡ2 [�j�b�����C����]������u"���`\o-bW�(ꛋ�Q��d��ò��Y���%$H�Td��Y8�?_��i��zI ����9q�s���3u^����I7��s��"
�Z�RHk���2R#>�4�&��s�x��|���B̫��Y=F���)l������lt���Z1'���wloiV��X�y�����M iz�c��>=ֵtw�h�N��V�G$�*���+
�罇�Y�ҽ�w�� �IUr���+��t!" 2��bQW����ܐ�g���%{D)�݁G{�u+%_>�5LH���K�6�C�P�0	�T�J㡞�4�Nlx�^:�I��8���O��� |
#S� DZ*�*e�����t���$��d٣��N���Jo��ڱm���>��������YM�F ~|%��]��l%R%co�PhQvPH>�PT|�����������d�]e�	�����}���6� F"؏`��V)�I��g9-w<�]�8|��.�`#�;#i���:M�}T䥹w ���N���
t
����@�	)OԘ���jHi�8���V����HlRR����`D�+��$l��1z��ў�_!�S���*�v�ݳB�#үsn�GY�=aQj�/Y�1�TBB�`�6lbbTߎ�Hb>]�(�1!? �\j������D�꬗C ���^�B*FHQ���}{�	p$� <V���ØW�Yz��?l-�ct��o-]W��|E����;���з��p���'����DQ	f��4�t�
�L0r2������~��q*����7��{VGGݣ��@��XS}�sY�'d�F_��_�� �*{BҾ@�ۂuZ���
1:��{���[�]�����F9��#���:��Ԕ�ׂ����6��r=�e!@��g���98)T��Dn�dJMA�퍘��Y�t�dc�W����g��K8�e~�&���F���A�,rl&��͊;F ��������b�
�P2�\�l"�����Q/9%%^��$�8��Mc������w�HSW0G��34��*��A�1]��=~�T�	4(�eqJ~J齰r��V-N�>z������T(�������E�ߩlήu�5E�{n��7M�+%��-�<j�Z���4�&��`Tb�1���A��m�R�g.$� ����N��eN����� �,9`�I� Ƽ�yyK�mizM�h�*]�T�=�� Daݒ=J �o]�%� �3�6Gк�JK#BZ����X� \�wO7����FQAz'��-wD�����ht:L~��0p��||�����A T�����+S��Ync���{�����q[V�*�s'@bTQa>e'&������qSH�`���}g 	�3;@M���Ke�/���%��g��By��lwy��o�-���<$�g��)�c�j�ULRC|��	ǅ$����5Bkrj�`�u�;�������*c��2�C;$�"��E��?����t6����spppi6�͖� ��J ��/d9_�(t�koo�uV�Xgӛ�er���}[�?�a��YF�(f��}�N/���͂�sV�{G`8�OW�5f��@�&��`�/<��|�:$$���r�3�]@�L7,��t���\�Yb�D�;���YVNnYg�8k�����bU��6�ؾ>i�4~U0*%%v�*
$�j���G J�
�YK���m�Jz�\V�8��<*,Ђ?>j�l�{~}��ď��F����VgR�*"���C���͹R�b+�q�u��5�k��Nc���t�B�~Cx%mJ4V�K�x4��R��5|v�oe�x|����:}P����,a��5��e�a���թ��L�b�P^�KokW�̳Q;-�U��f*���<�~pP�'��_����P�����?��8�A�N�:x����u�xZa��-�Z�j�_��*
����тR�ʛ7�����.�g��	��ZFqq���x�Ąr��!�#��P���̗��	���3��~SV[7�ӄ�)G���($���T�^�t��,Cq�I������JG��֍�n2$$$i99�C�iV�)���Z �rn�9���%}O����-Y�{���J�+sbA��M>u�����%��-�Q�ߔ DJ��z�(x���S�z^
�^�z������6�����:�N�������"$I�a�d�q��Ėw|u;�?�ȁ����5/�CE���|n�9����!��-.1���SݶM�����S�S����N�_���%O�~���|ܨ$~k�ޢ�E���h��0�n�?�n��`�ݠ��G�Z7j�͊8�L�X�
��?�G]�x(�T;|r����S���FR��ed�j�8�-	{���MD�4)�;7|�k�l28TSW7쏦v�H�g�}�}Ӱ��{ٌ�W�<TDϔ���7|c� H���κ�J��L�����K��R�� �P1b:�������&���(
����x�ٻ�,:�4�I�]%7�e�ij���F�I�����v:�pX��.%����7���}_A�pY۳t���`ab��c���x���	k�ё%P��
������.�Cּ �����?�<^����5m�9���e/����?:y9�O�}��L)�����޻�C���d6إ��W�C[6�v�����,��\�c���X�Ts�l��艉4Σ ���
�ǧ�ޅZ���P�j�mw;)lᰱ=R�
�/�.o��h��>?p��oh�����[�%��tyr�t����l�}M���_H���b�v���		� "Vh�?]�bo_'&��b 
WII���6���^��K�E�D�A�|�p�����)�����=����Ԏ�����Ƃ�k�a��xe�Y�|}��g:�5gP����d_���jp0�������_�s¬V���Ô��o�>��f^9Y���Vf�?�P�.�s�Dˢ�Mi�$:[�� �߽;@��������� �Ca�,�9���1x�7��R��0���w�gw��J���M405�Xb&��,zC�|Kf&�o�����\�m�ڢ����p ����Hpۑ���������L��JFp.��,��m������%'�O.�,�sq�h�.l63�޿o求<2���ʼ�h�`�h��g���=�G�M�~��q,��;+��vC���޿ }�)l~�KY~�Y(�S�UCD�D���-�}�)�h��#���fT�狌�oWm��ֳ�W{�mmR�fk�?��n��{�&re�a�(ً�����/@,���5j��̀��sޏ��`��V�C�������`{�5�r�z,��o�rs��q�q���z�W\�*�㪫�H����M(�R��R7?�ys�evjJ�P*��d*�UҀc�B���T�Z�/:����b��Rq&��n��ԏ H��!���{^����u	�����n:MM48|O6�g{�ρ��̳�a�5� u ���pޒu����|���{���YPXX,��R.@��uti���Ǧd��/�_�>|@���#-��Z\*�i���~l,�����ǀ�8��Y�s���?��,��k�PP�{�FJ$dii��;�.�N���.���n���<��~��������33k��ֽ�{�!S�2�oU@12I���?݅z�F�G8�_p�����t�����Ɔl�9��
��ZX �ˑ��E���� ��Ů(*	z5`� sf��
hr^��7`����P���!��_k�`������i�n�ԔU3�����=��������'�M����2�op��|���}��%���J���4��,��J�ʋ!?�����>s�tLE�M$?����Z�}h�o�߷��R��n��ڪ�K/+���ٯ�
��_�҅@���!��X+�d�ԃ`x�w3fUM�""�A�( ^���9N�?�Wm6��Pc�/�A��7TV��'�� ��-<2u�9P?��Ġ]%Џ���*��5=���X�vH�������3�I�����?ГrY�v@=a�����+I�1���!��fv�[�I�j�(-��6��Az��;�d� �a�׶�Bj�z���.F��? N��Љʭ}w��V:��m�j���G''sf�`0���w]LO{�i��Avۃ��"Vr1�����gˮ'�����D���Hd�%qYA�$0��47IIDn������3�W��i�"�L
�GGw Ԓ>�������c~ш��@>����RܰsC�v~���O��@4�G�\�]7� ��4}^3
�â�΍�ԢY:��%p��qա|�l�}�OtY�,��97�'�a����"*�t_�6l�|�>�X[[�E���B�C
l�[�%�٭�EE�f�%�	�2�g��\�|H * ��w�Ua�	q��K��=F^=H�łV���BZP�%�^9} ���t<Hz��9�хZT�dO���ljw��xj���%��t`��zL��2W ����{�7����64��(^�^G���v�� .V�|�y�J����ng�O�,�C�o��e���a��ʹ7`8Ή�yv�E���<�n���_Ťl{:ox�%���]o���@���?S))��0�Lx4򋋾1����K�)���3��XP-@o���^woB��Y��nhUJ�b�=��+ �*��SI���Xh�(t�-�?�}������؂K�:G�l�eq���']���Wэc���OI��m�,�x��7��K=�`��8��E�O�PN �nhj?Z�#s�3��4m��T�����Dҋ�Τ�cQ�Zpl�)�R߁�$���І�'�`Wjў`�V5�#{Uγ ��|	�m�|E.7
s�sg��Dh!�`.������ϖ� M ;���;�P�w��v�?��4��>����� ::�zFñbQ:��ԯ�!�Pfw]����/�t
=aLQ�����$�쬧y��Sv��W��DDK ?�wl�+��f�%dяYZ��֠3>k�r���Av�6�V`jw�����������_����T߿���k���hr� �`�h��.����Cw���З������T$�0���N���&�:nn����]�B�$Z� !((	�)@��7�z~�q�Rf��	f�9��5���Z} �ܔ�|	)�֏�d�?ήo^0�?ӘZ�ht�~�gH�A��Oo�K ��f�P0�$���Ia�9i��)�Ϛs5]ϛ�y��񾟟�]{�#>~ 𸁁@H:�������c!�￁���i0M��* ��C��d(�n� �a  g.�A)QQf;�t�W�z3>�����"�;ĺ͒����!s����)R��4O�O2�߮`����xS{{��8l}#$�@o���yi5��[��+D�U^��E������O���ӥ!�'-j���_G�mE��9�eu�Ѓ�FiH(#c4��NQAauJY���K���A�,2�T(BG��P����@�j�0�����2��.��G���4�T�\�d�Ȁ��,���iI*d��٨ͅ������u*�����K84�T�ї���<�Ma-�Yb�F����i�j/�?��[0�����.m}�̬� ~1H�@���A��{%{32��}�������,%iX5<�a��=Ƞ���� �v�8�b����� 
���Hc�33��رa�/.���X��!�{p�Z111>�2�M'�ە(Vb�t=�$�wQ �d$Ȼ&��ֻ�ʑ��X�����T�@u!!!9���"p�3�j�nw�Q�,�!D�yxlw�N���	-���;0M�{-g5�(����M�.��2ͯ�)!�H���Z{��*�t&����'i <�V�Yt9�J�q��SR�p"
��]Qӷ�)i��J�OS��fTm���� n��F�"J����=�t0S&�̧#a�dTU��1Ol�o�I;�ԣ���%1��f}I�ʄ��d �`Z��X�jP�Y�#A[����m[�By���o����I�߲]+�]� &�FÄY�?����� ���Eu�T�zd@l�ZZ�h�)�I��V�cc��}5��ь���hN���3��u�^�W����`R5	'9��;D�C���m1�tL\dz�)�KO���?*(����2�O�i�a:��ۤ�",��Ĭ��̢�`�Y�|�S���MEB�������-�N�k����%3V��<��fe�--��ͭ�����	}�]}�������x%A�Γ���C�z��2
��Zb�v�S;+G��m�0���.SA�y2����5�6�
��?����X;]����S�Dli~5����YDC#������>�
�w��{����;�/��Z���Z,�\�i�xj��$��l�N�a�h�%�j��9&8�V��s����# d�������T��+��@Y"V*�Kί��L��$������	f��S򅘖�����(M�j0��v9ˉ�}��sPp�?�ں�io}��We�ٸ$kfM�$V��jE`3�����S?��5��Y��ʎ$��bh���MNN����\/1��+�'<d���Ś����q������e������1�̍zY��h���;�&9�3z��o����A@����d�Jf���Pҥ��U����}K�<�},l0e���$2������;���g��I5� ]4T�w�c�
�����O� 9�ڪVR�~Yv�����5�.�R��ӫf��
/*��4���u*f3ʉ��/ň̢|��%����{��7�|��â��2�yڍT��̖����r�������F�Mv�z��v�d��M_�<�;���j�04R�@@	�4`ߖ��������Ne���Uk\b��� '''��n�!���f�J���C��l.�Y/?d��+�-V����{bb�
��9�]>��&���D���MU�2��c�<���=��D���P;SKKq%��CR�����~�ӹ���Ƙ���=�=���7�\�vǄA���->k�ޠ��l|J��bK=J�����)�9{�+.j&�,@i��3�2�q��W�g��p��[x�����[�a*�N���T�Iy��5�,�H0x����S�׿�|�X��7��%�^	2wߩ"��qS��!���f��+���xP�
���Z��b[��ͻ���=u/�Q�G)��9�ǲ�� Ts�(/��=� " w�CCC}}}���.�y��\�9v>q���'��D����'�S�l�F|�-V(q|h��My�E�"1��d��H�ٚN������`��H/�PR�g
e>�u�|a%�PGp�H�Y�k�!�ʓTѥ��:��s��Nw��$g�$���W�S�/Dc��1t��/E�d��A�z��{���)��+�$�)��w |z�?�8�|C�0�K�:3:�u{�C�ͭ��_ cs:�&@9v~�,,Ddg�s�N���.Pb�TT��MN��,��P�� n��jm��0^� �f�\��`RZ��bg�wBF�f��JN�,e���	���c {���A]�^GxAFp`�q~-<�SqC&�tu�CMDU���`�7*e�&�����Y�����$z�¨�K���VR�9�gF�e�Y����x���ZG&,������|�����'D����$�8ܾgJ\��Ŷ��;�Ȅ6Pd:l�V�*q���~���Ѡ�&�F��yvm�k����69�+yWPP�:���ٲ�d}� ���I�|5�pe4��]�Xd�x53~�Ǫ�"v��:'�ׯ�ng��u�Ǎ b��o~����,S�u�������7�mJ�*�w.:�;�?�9�]�߬w�Ձ`RX��,F��Z�t���wPyr��HM��3�tޟ�U��}�t@��G\!�u�["5�_T��y�as��A���V���L��WL�b_3I�uo�c*�m~�����(��'t�9����������L�?���۷o��V�KJ��_IƳ���X��$5LX��<j����VK[���8�� �A�U��p.(.~-.���B,j�G?~�=��m�V��"����}L�W����cUJ1;r҆���[!HL��8���-C��ž�NL�n�?���ֈ7xE٪�Qj�TW8"瞭�v�vL��z�e��IW�[�Ə���?4@��p�(V��=�|��L�����y$L����-p�Fi����<0^��nO�; a�P�]��M�m��fך��L�F��ѯ�d ��ܼ��ݧ-��LMMO�z�:�l�;��~���/&C!P �%�����h7B�ã!�L�<�ե����q��>9
���^����o	ލ̾��g�&.̂^��:�?�+vC��� �M��L�B	e(�����{��-y݆�5�����$�ܿ ���3s� ��k���� ������MJ5tQ��7�e���Q�q|�w�ޭ�:.��UN�\Z5B��A�}%S���G�+=��:�~�GU��B;n�~n��B�5�`���²Z�Ng�">iՙT���$p
S4v��ꋂ� �J
s^ ��v6�s�{����bXQ$1e)�'�����P�8_�BɁ�9�N1q��0�ZÁؗ�V}^yj���oߪ��A�]:Ɓ8�Θ	d��o��^����.ݍ�!�SH�wh�EU��YP_��Ύ�Z�����ZՒAO`�r�)��.�&��H�B�JFE�{�AS3�
%�zt�K���	,��Vɉ/�RF�$J�QDĎ58
�������!fe销�2�]�׼��J)n��u8���3g��ޫj��X��@��<��KyW��踱���-���r�\�����ZJ�oxD6�cu�7xS��\\�C�+]c��'_D7-�I����mgdf
]-ㅼ���n�AT<9*�$N����cV��Vl<�-r��wz�B�ķT*�Ŭ��%�F��o�XI||}��L+X��2wj��\Ep��) &�@qG^j_���f�YGn$ X\���Ϸl�y�'���eddT8p^�z���X]Z�(�p2�pBÌ�:��4�X� N��g�+�6��5_'�`�sw��c��k�ϟ:���@m�k�0�2���N'U)$���}��/ݛ8ә*�?0٪�0J�?�� �ڴC��(����g�gO�S�r��XB���G�]����=Z��E�c8|���1��C���7�l�S�t^� P��K�R��}USc*FǌJ�t'�|�\h�sҲ��U���k���	�z��G�(� 0CF��:��b)2+����W��}�c,�5՞����" ��@Iik��&n�Y`��ꮏ8iH���� ��(*Ieٶ���Q�2�"_>��qw#�,R6��*�ڍ�"��\m��R�Yi=C��7�ox��v�#������X���ES��!�z �Jxk��r���b?��x�w{�E�̬X̂��k�*�rp��ƹܟB&
�ͣ#�s��hO������s�㌣������l\>�+���C@>9�h�Hc��wS�|K���O:	�;���_V�a:#�(�4׃&�\HY��v�{zV�r��>��/5[�����B;�0j�T6��>���"?P�#���{Wz�za���X���5L#(HVi4"nk��'��~ߡ��z�j��=@��2�(�_���A�x�}m6z2=��؈�v �w��=�#�Yts	V�|�44kȬ��rZ��qԬ���\~z��<'Ñ�>��;�'������-˼�ڵ�0��F����;J��4�g>d!� E��RF���9�M��J!��D��5.Lz8�j)x2':) 	��&P���Z�sK�,ML_X�7w<-�jY���CҬ�t8�M{�%�?^ȯ����JNF����<��611ٝ����ɘy~*ba|\.��N"�����EiiQj-��]*����\%]�Á��~WW�ÈY���PU�Sx��%"�����UK��(�Y����l�Ȕ�Q^����QZZ����t�G�ʊ.Aڝ)�į�V~\<���'������ŧ�?��w��
�v���l9L�AL`�/'ť��Fs����������� ���}�Ⴣ���%����FG�}�}	
�w���(D| ֞Nc'��`Ӗ�Ce+>o�ͽ��z�����c3�-�&O�-����Gா�r�H����h��
,,�u�z�ʛ��2	�EZʻqqx�FFT`0q���hy9[��{������旔�M��w��R��(mnn���!�n��~}����{RDd~A�ڕ�דFNI�
!��2���saU��.Po֗�1fv�� �\0U�e�6$E���(�1[��}#|mw�!K�=P�^�|��h�M\�����&?n؁�#�5V��ĳ1� :!��`��%J��=���%- Y6A�(�#��^�m�:��� ��HНr��=QEE��`((�M�󰧦��KK�@�F��W5WB����׮�!��x��׺O7�6S/Sm:wq������O�j��ffh�&������찢����k,����� ��X�X*HE�N:���4�M�N�^ɞ0]��|I��^��.�͘�~�B��݁����-S�^9���p_�����'�́X�q�����Yw��c��3���@�(�y�חj.$��-Ɉ�"u�����/)�x�ma�#�Zu.D��/Uu87]� FF��oh�ު*yGW�@[T>��/*[��_��ͭ��5�C���0��fT:Qo�>b�Z�q���)ތ6��C ����l��ߐ�e�Mx,I4�4r����}�����W����.8�O�o҅�Bp�TD�,O�Qz��RBrȹ�}T���w$(���]�ݾ�LJ�Baj��\u;�N��6��^��-iW�=9'[k��6<�߯��ā|���;#��2ȷ�1�n���M"A�I��n����w%�=D��[V��P�B��Fo~.��8j��D�LJ�r.��O��P���}z\�`��u^eh���lnb?���܌o��iۤ�ju�N�Li��i8ٺ���)�%��Nz�+%z=�9���K�3����=c�_%ݴZE;�I� �ޔ?_v�m'��r���%(�As. �V�KI�_r�}�R_��7��*+����ɗN��Q��:���]R�ϓ���n_x��f�rc���{f��_(:H>kkL�ɪÃ�~g�{"$��A�t�Wऻϑ_f��G�<ޭ��A=�Ji[9�V%�����C���N�Z��q��h��W������Sdt9�d�g9M#LŤ���K*`�j�x���;�%s>k����PO�Zx/ x��)���2bɧ;��}Y�9����vp�Bn���(�o*��[�q|��Hfhު,��;����}�t|S`���n�H�|�$�N���g��$!^R/�:���;���O�ׄ~�D���Gvz���c*��YZ�]|�FHa){������xٳ�P�}�/^��H�I���mGk�=��
����A�+�%6�����;]�^rA�^�S�W ��Z9�=/^9O���s�����]`�>�����(xj�?K��'g��iW�vEuѰ��X��j��ymk�OO��h��ߠ߰�H��=�?��cz�s����u�Fwp�(�а�"'?E�� �gl��s�p��k6D�<]'�>��R�BY���m����w�v��^2Y�\�K�*V�lD��2Z���v�C���4Y��QV��M��#Ϫ���{.�z��C�~���p��{h$y~ؔ2�l�ȇ~ߠ�]�}�REj( B������֞���ʟ��������
J�e+T�P�;�q����)Ԟ��_�&&u{��,;Պ�;��V:�<j	�)���U�x��r v'�'�ɥ��A�P[v��3[��K�x%��+3>���I���oV+%0_F%�P�Nx]�)E��[����f�P|$ݽ����25������ b5/�C������3��=���^�8���pv{���!��9џbX;Q�5����{H[x�O�h������]~A�ax�'��,�WӔ�X�!���R~~�� ��q������)�!oi�N�W��}�������حN���xˠ$o���B�\x��k���}a���5n:����������� �"b��H�!k*�.��O�R�̈́�=Adʵk�:'���KY��O��77���9m��5�!�7�p��%⩏�:�}��U�X�{�k�/�J���C^�\��|��F�wY"�C6UP�H'�>���`ł����`�D��Fif�`Q��'������M�R������V�1�����V^4��隳R�έ0y[h�J������x龟͘�M+����S��87瓷�Ac^e��!���٥�>��
��
B�6�l$xle�Tc��
s�ސ�I�|T�A�qoY�̣���7��;:;O��R�p~�����ڂ�W7cG)3>j.�*���j��d�{�nS	 
=���y4�{4�mX�Xē�
G�X[�[TM�->8<.S���W�H�eWkҤEDZ鳻ϳ�Y$V%�00����Gv�z�-Y���;7E#��t!�
�T/��Sw��g��Ѧ.�Od�Gp����4�M��}mY��ǒ/��e/�?���8�k���^]���=��{G^���m;6�CL9�T���7dO�Љ�u�zr[��%t d��?faw;����7�{$e�J�	��*J|��L5^���9��6��;�z���Kψ\&|Fzt���^���J�b�#�?�ғ��땠�8�L׮P+a^$��vH��_}��p5�;�O��e>�;��jr�~H/���CD$8�/q�Ű��h �M~�i�1E5�o�*[�y�Έ�=Xs`�K�[���Db�Px��3�a�QKh-��ՇX�KN�h��M����\�]Ǽ�� ����UK���xQ�7_�aɔ���s�J���zf���Ҵ?N}�-��w��	��K��N ��̮`q��f�U��������m�{�;)�H�ZC

��M$�N�l�6�ts"bc]�۱�#0ߧ�Vg��g5�G_���<{}YB����LҺ����_.m�����
������zM���h�;ewGʘ�קq�M	GR$�\���L [�\��W7�����W�̷ӡi�5w���@�`���T�*k��O��x�Kv��{�]{K�e�RRϦ��5%�͡�f����H$L@���czǇ�ڴ=:�KVa����k�kFy����M��,f�Ʈ����9�xht�tr5�@�oa��,Q6����E���탉9#�K-a�1>j-`�I�;&�ӆ���_���h���pbxi?�sB��,�t
�{�b��ٌ�9IGu�bX�T�	9]����Z
S�@y�?��VJ߽�RF.��4�����$/�&�;M�s}ynօK�w�;|Qjjᓨ�h���<A�s��Z�@9�w���h�������z�m��9�PA�p(�f[��U9���H1U����}�]֌�X��,AXtL��Qm�Su&�T��LJ�뉥}���Is<u�61��J�$+�`�k��ɘ��ί`>9�IT&�K��7�N�����,�D�/#{K�ŀ_`�O$���4�?gL͂+���uy�\�h����k��W~g��^�gEH�.�}H���o�B�l��3���W���q@�G~*�eV#�����l;3�L�Y3Jz�ЖM�㕯�w:@s?�N���&ҋR�Fe�Z�c�1�mk��*�n&\M��/a	S�MՂ��0�t�o��`o��ef^�M�b�z|
(nBlz%U(�4�^�EE���?��̳���\��ݞ��8��^35��g�t.pwջ&.��{�c q�	P���wtvw!�AAqP���h�	|���HX5��N :zùݠ���?��S p�zy�EY�/�; T89R"�v�fw9��%������ڴ��K랼��*[dI�����/�l�e��Ţ��~~��}b����鉚�҉_^��x��l�(���Ǩ��ax�L���F�oZ�������Ez4A���Lʇ��k��*b�=ӲOw<�]�2� ��qd�}�j��տ�`�ѧy��W����#�� m~�1�/�,��F�uMħO��d����D�(M���{��eO�'�G1jZ���"��.9(���L��OeAH�j��9���R&�p�'v=�#�{AyI,@��0��E3	��p���pa��R2�G˟�
��"��Y�&8�![��Í�$&��Ѡ׸z��b�Z��dF�=�yn�������B� ��N���Ah�bGoz�O��EZӖ��̻�!vg��5��h}ٌ����8� �^�֞�xu���oŐ��Be�����)]g��C���(#��8�6®�g�v	@�4>�E�Cz�:ڶ��n����v�0��ᇜV3]��~I��uD�l���E5�r8�����)�1���� {�Ӌ;"ql��o�xi��(���K:�"{?��7��?R�UӗZbͭ7�-y�O/X�){^�҈s��gƙ��s��y�0Zn'�]��#B2MþH��=�K�Jի�B1���UDS�t�]Z��h�>�n� I��cʒ��	�,2��؁��q����h�h�����1����wF0[^0u��NZYE_���Z���.+�63G�ζMc���X��V��s�o*���̈���_��{Jyb&s[v�3+�8�HZ(c��y	@����0ڷ��v�`�(?by�Lqy\������3��!t������	���g��`��7���t ��������|O�Q���h�<��$�R��~���mSPg��Jp����aNG�:*���$��ށ�k�<6��)���Y�8�Ys㡹��4W77>���RR(X��P�srhE�0�&��pX∇��p���g��*A�DD�3��Qw�D@'�����uJ�*(���"��?_r%����===�z�Z�M�;2..����Y4M� �-o=b(w���f��Lե}��
�9O�Y�HH�-l2z�N���·�9C������9�7�G?���o�.Ś񜹔�$\�vɥ�dH)��o�'��A%jo���k�z`Rsn|�N��϶���Ő]�3��?��aN��y~�1657��!�"~��I�7�����J_�r���Ro��
;iU��])װH=T�d��$�YqbF@�gg}��\���9Z��>�Қw����?�^�n��q�i����+�vΐB�1��%zwۼ�<5N��i7e�5Ӝ�n�"_E�_���;kT���1#.®�rg����� l'�H�^L���a�5X��o�v�C�Ӛ����ȼk-A͘x���#��O3-��[�HQ�+�A+R� �y����(ճ��4:��<\���w�_�7+�`�^��d�-)��[�4�` �c���.}���?%��}[�P�~�F�F�. �]:1�I����[�j4/�z!���eB���fJ�0��͜�?Ӛ9-�#$d͉ 6�.��>>s�&cN^@��PFd��lR�8��<aY9�㮬Ŧ��+P܊�>-䵥���y�X���
Z�@MzWC�_�A4i���K���R�1ܫ!��f������bf�7�.Jew���Jbf�U*�G.�*�����̞-�)2)��#��f�%�7��u��=tcV�jDF^s�}�<�Jā�M�ܕ#:g���0���u�j3�O�	�#���r{��Z��2p��u�b�W/2��pR�vɨD伪�n�E���>�����^���%��5��I�Vr��B���Q��	k�!O��";�F���ժx�N��r)�ޭ6����2��w����B����HB�0�2{���NG����s��i�3���m��ϡ5k��>�g=�V�j�jU">O�5�A�?\�u{���b��&󏟞ꡯ�D�tj7�/0�!/�����_5E�]k1����l�n]*Ux
~ئA]�R��$�s"�$�!�ka}�Qk����Y�Ue̐���p|�>�X�i�,z��l���7l�'c*[�
�ܟ��>�vv�h���8!�B�{S�i��+`���=Q���R�����R2_�[E(14բ�cΛ��b�.�o�S��(��ļXN���6�t�v�������3
�n-��f	U��p��|�>q��� y'FCK��է�����A/fV�)�a�5/r��Q#�+Y��9��!,
ɤ�Բ�/�t�d	Gi&K�=�J�x��V�6�/}%&��C_a���8�"���גZ**E�;+�r
���ό<� G���׍�oBY���^2�R���Yg��Be�Z����8���o�]�[�{Q�99�u�phi�o�#n,;+�I,���!"^���7j��^���>A��9:3���*k�1��m8���e{}�\l�vԷ跾��/����6n�1e:������ ǥ`��]�i�M��'����Am����]�r2��Y��g��c��$vD%o:����;���s���p5�-�x&9�>�^�0�/ΰI���F&U��{Y�8u����~���d t�i@p����z�Ms����C�����^���[�O��jekK��xKF'�)o�0�r5] �g>�/�J�Y6�K���Qܯ4>�1��/�O|��$�������Hӏ���$��*�e�f�?�h�]�f�
9�1�,�a��S0�C���LE�*]-C�ޙD�8f�RB<�>
/�{��mr�fݩ��j>{՞"���d\�c��nƴzw���z�[ͪ�����ZGA42��T�U9
����=�ݤŗ&&�K��.Wǰ1�w�b+^Z5߆�=����<�8T;�]]'/h��d�����s�ߟѢF]���&~',^�AW��_�Y�|���؟��Ţ301���GT�j+��9`�d��e?��6k)kiѣ��ђ����'�G�to��A���n�2���K�xQ�uT��N��l~k��-#ˌ*��6�D7���3��H�҇���ˈ�hi�4U����f!�e-|�������A;�OX�#N��Q�܇���ڬ�]�����j��%�w!���^�܃����(.&a����L�	�]��M���ԧΣ��[8��z�����y�z}��[�4�$(���ξm����J� �a�x���/L��d�=��t@�0���EK1�r��RpF�Cf�����	�N��C+���?�zH~�T���6�����cfg5n��g�m�|ޠz�d���	7�x+KT��C���c�Y�:Qt�;�<l-W�D8Ih�����4?oc*��s�d��9��Ҭ����G�ٰB嫪���_����M�$?p��ʞ����z�<�����`z	�BB����C��{w7?�9$L\]�M�jEH_{U/��v�%��SH>��L�+J��/�&k��0l��ۥs!\���]#Y���7\��������t�	|��Ǯ�AFJ^%�P�.�I���8T�	wB�f�<=k������4�3e�߬E�Z˿�8�����W��8l���������fc�Z*��d�o��%$��WV�R�wXR�ogL�9D�ѐ6�D/�!
B;C����r'�R�"$�٤�}��َ?] �T��Vs���z䨀���]�؊���9?.�jQ��W��EoJ��;aG��o`J��ѵ̺��Єo�׬3�Y(|G�]��$����5��z�&BeO��BV �4�N7*���I*��Mޗ� j��I��yvH�SeaF���<ԙ������X��Ao��!K��z��̬,9H��~��k����
�[ֵm�Ww�ןʪ�Eg�VBmPo��yJ��Ą�ς��'��ɂ)��z\����Y�|�X�gլ��0��6����>bv`r�����UF�h,�/���ي�ٸ~/H�T+|6���ˠ�3������c��w�8#Y�3�pne��n���7t/]�곍��8�Ju
e���Uc�T�f����#��ڂ�PNǳ�Oz��+��e�ŋ������rB�XO�n�ؚ��D���y����<bv�.��l� ?��I"��YׁH��=:*�3�ߨt�M�5�e�;?���}��&Z�Ǽ�G��[�|����i��QE��ϩ��A�q�U|�0���@Tؽx\�H(�{7��l���5��.��q4It�	������ov�]�.-��Y#zⱏY�hJ��ɋ�s�*�q�c]�J:��V�h�|�J��l������-Y����L_h���rm-x�*�Y�Z�@3�ڹ;BzVeYԱ��FR���O��;ǭZ~�|>�/���u�K�1ԏ����i~�x��]0��Y��d"�r�^���B���9�B�8S�ӤW#P�����<wN�ҟ��MQ?%ty�.1��.Z��S�7�9U�Jḇc�?VC����~�nu�n��j-,'g5`Wb��i_��9	��¢E�q����`��d�K����)���ۨ��Q�烴bR��%���	v>�0M|���l�>�H['�"����9o��͆K��y{a�I�t$��\��ǰ���-0�W��|%���н��z n�)W�H�r1)�fѠ�&��_ J��pG��uK��<?�h�������W1��	�\�J�嘻�-�Y"�d��p�ĠJ���B0|�٤iA10�/�":M�%�a{n$�nR��_R0������
N,Vj�gX������MW(���}��S$!���2٠�Ǌ��y�Z��^�e9�,�h�XNȂ����_"0�o�h�Ȳ��x����T�*"7�8��'��.B���z(�F�Q=���f\�e��s�B*�M���5���l	C�B#D����O��T�J�1��[�ߖf=}��U5G��OD!}o(�y]c�@eq���{QFR��pڃ����o@Ѳ�0
\h�k=�N� o��ڤ�+o���~���'��l.̲��&_&o��0�C_T�?-���� dȹ���kI�\Ό���^w�y�\u���f������<b�}�n;iō��«�7˲���j.���hV��^Z!^�bA�Khd|(�`��΀�����1���UNi{&G�um�0��Pf���}���@��<��]��t}��"��U�2#�⒔�	)x�ұ�͵[�G����O����1���+���?���h��x�5#�,�1�{���M��+���~��X@M����o/�O�]���Ц��ݮ �ǋ ���g� �J/��ٮ]�Б����^�����+�KE�������'�Z꾕�y�" ������z� ����[���o:R�!ґ1�hż`PV����u�6�@�|����:����T���7����"�)2��mK�h���O���v�n�o`3�<|G�x�IZ����>8��P�k�A��ۜ�F��Q����X1uF��# �lʼ�'�ȤO��;m��t!�L�D���٦zw"'���s^9�S|�0�8S ß0���k�m%ś�!�+���2(��0S��%fq����Lԅڈ��x2)I�����sT-��Π����K�}6��f'%�W)�a{�CjGOA�X���3E�E�K������|mK��[4����4ys2e��_ǿ�d�4g�j�y��w~���d+tyu��^ �Z��~��;J����EA���`����(��'MM+֊�?����đ�Ԥ �9'�����U��-Bc�_<މO��ru	]�g��KǬ�R�͸`#)�I���e�NÀ� �x���[���@$��W�1��4uOt�*E��/ެ��p9fo���Bz7�:@3�i��$<+?�����!{L[aĩ����Ϗ`�V5�����t��m�Z`�;�S�=�gm���
��W��bf%�f�/V.%ة�6��j��W-�%x�2u&&���.���W0/`�l� ����l��%t�QW)r��l�� ���  �N��`�\��o!O"{�d�.0d\F&J���h��G�`q��0D�3������:rZR��/�1U�_H.�>�:�۫2[6�}�p�8�-}�^\���i��|^�{��#u�p�o�Ca���A�d�{�:�)����LOe?���rL�Y*�r^tv5-_x��m���������xe��ƚ�_f���7'c��pv﯑��O�_`x#$��1�%�r�<t����Գ����l�!�Q� K՛��J6d��G�^]���a>&�3��"�4�NSZ�ȾJ��R*z����\� \��sy���g�`�оh��N����!��[{�ֺ,o�Ny��2�v��À�=~	i�FmEwd�odh�$*�C�"J��o�Z9J�`�I�Q��(aBtT�����ߵ��?{�j66��7�{�k3
������. @�.-��� x/M����cIsζ�U�s����Ŵ�mZ��OO��0M'��a��`M��Ɣ��:6ύ.��Lx����a��=�J���)*%�ʿ�{I(�3�CL��Ї=�ҫe�qA권f[�q��V�����G��������u�Q=W"r����f����}�7n��P�eK��6��J+��a��W	}8��L��\wNݭEÂp>�U�"K��W�t�-$�nX[�u.��(:ff�9Y��/eY5�|�=�Ed?J��CL�L����c��}'>�aa?5���g,�|��l�\��o������
�VUM�&K貉�6'��I}�+���������>5b��-
���4���}`��a8��Eřv�૿cOS$oJW����F�]V��i�:��ڶ5�AET�TP����	(�kh�B�:(R�H'���{G�� @BGz�^/�{ǹz���~�5�#Y�k�o�=�7�\{�A����I�rP��C��%���׼;����O濶o|��޼)��ѹANv��ɬ�_�s��]�۷��9�/��[9K2�]v�(����t�s	u������	���ls߮ݲ�Br6����z�� &��G�P��X>Z��Q��ʹX�mlHi|zC*�䋙J^���
t�|��#?& <^�a��T�q��V��g�&�ᱼp�k]�M����q�2$.�ugD��Ƈ�%�\��m�-�F�$ː�b���2�%&�cm� ��	�ݻ& %y/���?�L�����D��e2��yR>Z����K�q�W��%ߎX�蕧6���Q/�����G���tNwxJ%���Q��W`u�94W@�y?��r�@�j4��
]X�/��@��m�����'+��!o�6#xP2ux�O���rƧ���������ɽU3�W^�g.�_w�����o�Jez�$�tl#b�O�����%����Pzm�VW^����'��N=��X�������Jߒ$��$oF_�{�Hv������A2֭�X���ziBE���h�tha2�V�u�$����%�b?6tN=�&��)��|�tl���^�,*@ccI����J�x�+x@L�<u�V�ܙSUո_�o�����;w��Ü��2D�}lJj+V[e�M\t��(��> ���b�&C1M���N}@0�ԋ�e=�$���k��_`X,�B�+�=M~8��r��nv,��?�����~uZ�d��]ZWɎI���~u2�tU�E�đ}�'A��y�r�
m��>�1ڡ��M����{�Ku�o�����	�#�����G��� Ţ�������	>�濶]�bΎc_i&�^߬ՙ�i6=t�Q?dw[	�N��4��q&�S��2l/`�Wԯ:}�t����rh�[\Em�^~�T1��)��K��?<�i30�^�z�,(t}w&�VkK������T���
�O�S	zΞ@�~\šI*[�|�nЎm���#
VE]��(GF0�H�'�����rU��g���=��uH�Ky�Ö"�aK�d��ZVSr%`I":e�~������XU�C�3����Cdxr5��[��U/L�h�d��dQ��w��)�|�9]�;[-I�?W*gmf��^!*���2l���>2���(���b���k����0���ܹ����q���h���������#��gێd8�(�q�|ÛF=�ߜ�۞hS���"̥����k��e���q 7Z�����**7�:��� C��T��S��}����!a���1�#>L#��'*�?b��!�m�9Ф}�; n:\Ȧ�[M�eB�a��"a�?��T��Ƞn�ı��-��J�9���䎌�p���_�U�ra�����f��`��:�9�RY��ˤ�� i'LD�q|!<�� _a�̒��NV4��	��q}�����1	� ��p�x��7�����6{�32�J�ڦn2�@��S��5�sIٮ�+�OX�9�,p�=���G,y��8��4�&���/4����4�|�͵,�b��"��|�%U��d�e���07���O i���X�M&��
q��9k�ih⼓�=�'_O�<�#٧jpU�j�]}�Fj z D"�6���>ߡەJ�0���ۺ�h��|�桿'����h�e:�v鶼�o�;�r��h_����;�iz�Y߶�EӰ��Ҵۼ��4�#��XrK �.��`�����z׃��P]��V���o/�Y�r˚,V��������&ӱd���	��!|\{���
MUn�5��� i��cK%�rB�si>��|Q�[�M�VV��, �B�!I�b>�^2֘�\?��>8�cG���]1��Ku\ܮ�O�����ۀ�r�����o>k#2���p��ZqnHG���J��|H��'+�t�iS�m\i(�n{=�!H"����P, !!!�u"gs)������(�>A��ܗ�4�>���n���o��i{��?�	l,�~�e#�3
V\�|�|���	����?�8Tϣp�,l���|��}�J�=��E�Iw���![���������w�Y��6j��W��kW���'�Y�`;^��gyy���Z{z�{!��%t'�k>]�P����H�ߏM�1�����T�}�������E
�o��et\"���ٍ�R�sNe�j��aK���lN��#ܹZ�C�;��� ���;���	g#�u.�Wծ?��'\�g�L!�	例?������+�a]]�1ZQ�m�j���\�Voۢl\m��K��,7�
ԉ�W��^����NP/���ߤd����������5q��K�mW����,�`���9�+v��8�~�GË'��l��zȔ����i%]>���R�Jc,��J�v��f�ߢ���/b*?���:圃����1�����&^v�5��4��7H��:$rCg"2h�������a�H4o�4��mO�|Y�SƋ���\�~��m.������s�$��s�4Q�k�T��{�-�����8�r�� ���],dcFQ�����L�N�Mb�@��f�LW+�i�rc�{����,�E����
�(�at�s~��`�`��f b�0 �¼�y�Q���(SR I�>i��B=��p돀3�jS�\��x2 ��<�X���x������D��BS�,��,> �Ft�m�|�?�����m5e�T�MՍ��n�T���_��u���L��]��̓������b_�ZYxw�s� ^�6{�Ҫ�"�A<��h|��D#Vw��y���|
x]��䵬yms1cJf��S���y��f��H���~g���O����e�t�sģ �R�O�"�	��h��w. ���|���YN�[��kX�"YSeW�C��Nɟ��B�o��Y�Ͽ2SP�7���MH^�<Q9�
pI�̂&B�ø�L��D��� ˊ�=#�����Le�mJ$5�ù��h��������J�C�����	y�ľ�/�VbUZ@\�4u1�&��F��Xػ;b����HMd7?z\s�����=`[-_1���2��v������U�Ϭ�ע�|L����ǽ�h�#ge�������O{�vV��|��7p�j�yʇS�V�-2��w|���I�4�Uy�7M��B�8 ���&�_kv�R�@�vS�as���}�s&Wd<�i�.R�`_7UuF�8�ʾa�'%1�K}�����3lbS���~��9f��5�ZNd���P˧oR=�!�{��	 \�OKD��vi��2���-4�{�X�է�q�����|Lv-��Mi/�W��y(����x ��Ch�z�)��EK��J~V�*Ag]�ɨ������FUËMh� �k��Nն��קE��O��'��;2�ދf���}L��<z�>�_�'*4JGW�"|h���4ګK��|�.��՚�_�WmHUBa����/���49G:U	�ϯ�|�
&HƬ:tb,�\d����<#p3�3^��`���S{��d�	y6<�QS���y��Νw4��}Zg7vʑE`�	 ��!��U�ۺஅ�q�^5��/��B��|aO��+�?r�="CZ�a�J���)�d�0��Q����B5���hrN֝�Ť��I4r�$2��2btP��z]y���� a#�k�`�fYc���)�e�Q���(� �����d�>i[��v�V�m�Pi��-���ϟ������+3����3�/�v#g�d�������Wm'L��H�a��YRm�{��fj����lël�H�O&�˾صj�lu�DD;��_�5�N9o7�1q��FB�ţi�w�>�i4rZC��"N���#�f���:��)�c�m ���*9s�-��_Ea% ����Rǫ�r]E:Ss�z����%�K�΄���W�V?�)J�Ə����q��ow�!����4j�i�|PO�ux��!��0u�k0G��W�%�ע/ݗ��X�O��\-���2=1��k��ҁ����֗y��n�or�wM�bKQ���?��a�/1?�\v�1Kg�3�����l�;[�����fq$�}o���4��rm��k�*�*_;D|`̷�۸����1�~��MQ�WB�rpb�Y�)���� e�]���v.=f�sek���+0?�ZԊ��Z	����������H�u\r@�V�M�/������J�>�#hƐ۟w�&n�JD�c,W��5�YS>2(;��D�|�@{��PԶԦrR­��;�1Cf��[�I|�����;�Ǟ��1�ف٥����b�^"��N���u��
SW�����T�fJu{��A�b�:u�l����H�#�ol�~clD��	�NFa�ۈ�§��9��eO��W�Y��i#���s����s>td%L5j�b.�-�?+яPUn<Vc'\� x���aP{ٗ��J���Mf�[�p4�^e�U����l�R��!���n�,W�����d�������Y=1�Kb�u([�ː{Ӓ�f�lly���JFu69PX}�C�X�>?e���|9��%\�[�na���rY�N�/ߔ��N�Y���PͪD��ee������c��������g���$��>�x�G69J�/9���K����K�F�hF��O�NϦ�}s1�$�i�J6o��p/ɤ��N�lG{IKd�=�m��m��zZ���M5M5����ke�bpͅJq���JN�k�a�4ut�
-p�~:{��-��67k�̓~9���YOhz�4��@��t[��*���e�@T' S��6<F5��@\@+3��Fs\����T�NKix��r���Y4��k@�c)aa����Ϧ��t5��hY�i-'KḪJ�$��$ۍ�sn�O̪�庶m@ �?M]�E[	�|�������\�H^vJ��;��s[��h�(w-M�$ϩ�-"��R��.%�M<)V�okd�R����Y�ϱ@��h�ST2�땻������j�PZ�I��ˈ s�E-r���8�.�bW��k{��LDl5�A�t�#h5h����F�	%Xڵ8]���Z;�2�폋I�TD�| n܎a�4�l£*2��rvbF��~�ڡi��MJ��8���Q)���Se���6n2��O�xo������N~�Uh�U�HIL���@�_�ߎm
X�y��H*c�W���9+�W� ߀Z�/��J�)Z�W^�Sv_��}8��=쌔�=���;�,�\אN#Kx^`�LuMM��X����1G�4{dwfw 5�mѫ�x�Wd�c�����Wi"F9==���Y5M�r^��R���9��Y|_~�m8��bw���a{:����l�,m�+�}�r��HB�ʗ	��+�eOU�7&��~8�c)���ʬ�s�t�7�����x� �y� ��13	v3�7J��ر6��E���6π���/�k	⍁�pvW��pɍ��ޞ�bA'��$kƃ�Puˣ��*<oU���0��`���I������H��g�;%�(.�8s�X����dK�E��39/9^1��'ץ���fR?3�h�2���hw��T�ҽZ�I���LOe|O�D���T<�`o�SA��d��3#�r͉�b#"pâ�"Lq��ql��;n���y�"��/hz�|&@�7�-ʺq����;��E����[��%�Y[���Q�6g�!؀e�� ��$��*0�_�C�[��^�/�w�G�l�J*7�5�m�sIt?�27b�S���F��B�������D2�_��0F����`��n*˭��Xr̍�����@o>̖
;�C���:I�1��OI�k{�� l�ם�o�C(m|6�!����mS:�Χ%S�zNdg�=��֯j1�0��_�`�#�S�5�y��7��
��xWzE�証!hz�QJ����X�����;<�f}W�I�k����Y+��;��yV��T~G����:V�ީ����ű0���Բ�Y_�����n�"#��4�����=��gk:��a����G]H�+`8@��A�Y�+3o޿)�+���e3��t`ir��M�6�î(�mU��� b�îg�X�T˪4%� ���8�����qN�ĳ;��#^)�ӛ�Jrn����s��)QeYjNLK� ��λ������)��7{R_7e�A�G��8�pq�����5����Q8�r�fZ�^�*�q�d ^[cFy�k)��hK7���s�
�5�r�S��r������5�?vbs��J�􏱙�D_ҁ�vL���)�E��������yd#8��u��ƠH�ïx��X��G�lu�B�\0O�{����G�+��Z�Ŧ[��x*jX��>/���&��m�%`靗�����8�=Z�t�"� CK��T �μ�&�[���DU�h-��<��:\�;���(���"�B:O����[��u�����M��}�p��J&8(�B��Oi�)Ցl�H���AP9@���QK�2C[E��S0�YG�v[|Ǧ�$֬6L���E�,�&����������#"�;
YcSD%VH��8��,�W�W���-��#�j�^�ۿ��M�!-|�g��G�Ѹ��}ts�:6j���:��Ie������.;�#��D�(��6L1�͍�t����E,���6��E`av���5�^(�lE��=���p*u߆d�1�����؀���x�5Bs(�6*B	��e�r"���A�zr�z�2@�T4(P}���������B�݆�[�Q(�> �e�}��f۟w�;���¬cF#U�H0��>�=���TZ���H�H�Y��Ta��dz�5�t-�/!]��<Ѝ5��Cs���H�l���<���UN�ѱK�H�S]"_����  �WV}s�"�v"�X��?��;J���:��I��|ɴ��)��L_t��ӡhi�#+�m�6~{���Z�D.�DS�{ҋG�������y�Z�u5�hظ�]�.�5�����E�mY��$��:�!���̯UC+y{�
]"�N��6����*lz.������ݳ���bn�߆ږ>�5*H~��w/c���?]���2��+�q:�X����3"m(�p􎏹��v�X�L`t$q�)I�X��]`qx%^��-����M�uo�4�q�D2�{a��l�Ǝz,�.V��9!�3Աk�̵�����&f��f�ƅ�����m�7q�{�Nry�S���$�96C��); �c�\�e��/&
Ӓ�}�*�re� v���ۆ�8���6���9
S��E8�����:蟏��C܍:F�[�;���>Xn�Ї�,�B�H�{S�e���#67�� ��Yz"����&���~w�@�X��D5Z�P��D�bS;{����x�dlԋ���w�q�*����ؤ�%G��C��˜#�g�,����l|���϶�O����٘�G#���Y5�%����8s�-�yH2��~?ݻ}�>gi�'�x�8���A�HM3(��b���`Ј��9��?��QЯ}��0>Q�J5�'��8���vΑ�!-oe��K\�wR��}z�\�W<��f
I�5� ﺨ�ɉ���?���U��U���}z�&UX[Q����Q�i��[���V�C<7a:lJ��~9IB�%��$�a$��gӻ{�������ע����'b�H8P1���o�����ط��/�Gh��s��f������Սc;���L����r�
R%o��PK   .{�Xo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   .{�Xv��� f~ /   images/4d249bba-3190-4770-b321-fb8fc027a237.pngl�	XS��=��-��P��(We�@�U���2)a�)2�\�N�'"��@9P0̓��0V� �� B � ��oZ�����<}�޳�~ǵֻω׎�Yl�z��[1��9HH�TKHl	�,�䧙�g�|�+��f�O�f�����ly:TBB�9�練�'�*�9��F8�-A t��C=�{���f��A�ۡ����辱Â����{N���N������-Ү�7�g���װ��6���������7!AAQ�}�C�����w4����K_��������R�{�����j1���}{k�<��=1�VF^x�/8o��P�p�[L,��^Fi���0UX�����W�C�ʰ�e9�N��'�"�1����J3�����B���Y���@�ڌ6Fն|/e���YMFb���7Q��yp2&�(�0�6��j����Հ���_ڟF�Ǡ�����c�t��ZD<$����}��p=�bu�l1|�m�)L�N�Z�ش=�Qm_}* �5�)�6�dK�.�
�}s[\�g���L�
Gwj��Yb�>�T�n"X����m�Er�$	F6��fw�oV�`r�������AU��b9��X��E;Y�{��x�nް�m��C�qF��p�8ƽWW��^�tO{���1����?
�1�*b�~��wң�(VN�[���i{������ ��91��\�-~�sA8�O
���R�x��BL�ġGgº���j�� <��qx�V�{沴1��tfo��qҀ�aHW��@p��H��׳����*x�
&Έ��X2����]��;_�O6���P�Z��D_;j�g�9f�몫�fQ�̩��22s��ܾ`_�?���0H;�Y�\�ЮB� W�?G<�-
�ѫ�С'�$K�<�lɠ'�����D^��@�P>�p��9۸�妡��(�n�O^hb�^�a��:�*��GA�0~���A�̨��r/����
� ��T���R�>�z�
��2��7G�jL(�PL-y���J�#ݖ0|6\�ѝɒL
��/�=����FZT�GA�`���[�8-���P����B(���0��+:���%��<XǞ��F��ʤ֜�����t+�&<у�R��(l8r�9��~�[���@r��2�4Qs[������^J�+��s�
P�L�|�H�$t����Gl�5wZ���v�]7�௠�2����'��|n��K�NcB�������œ�=�O��7x��̹v	]�+��6�ryS���i(f�=a!Yx��b�;�퀖3Qk:�����m
c��AV��/gG�,��WQ�e��^
(��WupA,��}F�o��5�()�75�t��r�U�eo<I<�s7/��a؍;:�-�J��c&��>��:� �H�ys��q�5�oO��Q�E�1�h��h��~���p���/Lg48'�����yb��J���;�70�����Є�8�)��G"w�\���*��á�|<�1��Oq���5N�7��3N�	M�	�x��wJA�I�AS�_{�ǰX�4f"&-�nӒ��Wh7q�>�\,�z?�Ҍ���:�
���M({,\���-��\���ip������R+np�4ބ��������
��(�Tj	O�D��0���.FAÖ!X| ��(|�cA/x¸�bt(7��$v�'@���d� IܑUYZ�<E�F׬|�5~_�j��l�$��p��l L2�$��M���U�#܇�Z l;O�aV�\�e�p��8v�*.�-ʜO�%�t	��bA�3M��s7A=�	*e�&*�d��c��P�s�4��w � ZJ���2p�$v��ʵ/�'��QP�N���y�r�S�$��6�(�{��)�Ѣ|�1 ��"ju�౓؆�)��q��	��!�fd<>�B,�#5{�'��}S�;��d���B�x��~*���۲4�*��%�ݟ��0puEb-�����}����,!Ḡ���3jA�X@�{��9ǰkA��_u���C���Uv������8����^b��`���Z[{{NFN�����fR��M��A"
<p��O�̬Q���@7g�C����L*/���g�Ν;o���<�x���ӧޣ������fM�7�.w��$��x�p�G���e�\i�T��=��-��L����Km��*���'��m��t��Nc-�O���0V"���&����������Wd�nl����j/�~�����Y 02�s��]*����E?�'CY:ї�)�//'�������K*舃��mɮu3팆�t9��\R1Qy�nv󐁢�*p{�>���=J:��a�o�S�ʽ(���#0.� �-�����F��赶�֯i\L��h6���Nt*�*#3��H��ȵ���>F]PLla��a���㞞}u�#M��ȸ������ᄞ�R5^���[<���ZҴ�Uߕ{wt��dge��v;��� �ȋ�/5�LO���I���ynO@{?�.�,�A~6u0G|�a��P�=q��P9h
ix�~��|/uf�Jls����p�%���XGz�ٯ�8��Og��C�ePG�*ãQ/8��z���0�C��>��7��6Ӏ�97>��&���%�j(q�A`L��<	k��L1]`�����}=�R g}yᖸ��J�=��� i�A�탢��^#{ל�-h@��)7�2�K��W�^e�K�ڔC;�@Q��	ۤ��1����+�NJ�ݎ�yL\>Azس�Z5��k��@z�H� d�,.x=���Q^iS!�F���ȕ����4Ǌ��:xB8�Y��&�&��Zԍ�۲I-)櫋�����<6��
�6�i��W܍��yF��/�N�^TF������=�i��t��|`F�$˟Z�Sf@��t�XY>	*n(lچ�Z*,��C�k`�=�E"L��{6[����S��
B[�~e�*�w���`O�6=�8t�!Sq�����^}������fO��"�I���ΈuHޟͱ�Ep�mS:�#��d�F}|h
��V��o�/�SOF����8���$>���Q���l��N��3#f)'��rCe�9�Q-��s馧`���)&ô㜾�tHE37����wS[�&*�cJm�x�MY��}�cl��7�E�����b�A"]�.��^!��f��d�d�����Qը�2nz{e���-��w�`�s$z�%���E>�qP�w��y����d����`V^�Y�D���œ����˙i����| 7�yy�"h�H0��_
���숙����r�C. X�誀3��$�6Ͼ����R�i�ho�c��m��ZsKQj��I�4T\�$Pv�ހJ�C�r�jζ%��7p�C�<���.�㥧H���f ��AT"��`~�ސ�O�,��Pw����[��6��ͣ�
��(GnW9b�����T_���}�=�������b�� ���ct��2jؒ�����U�cDW�pC����$���c�A�[���ױh7���ⁿ���|k��4�&܄�@y�,��s�*w~�_(+�X�1x��$	~��=�u��aXL���F��;��j��&�I;�oj��ωf�D����\�3U#h��S�s7ܗ?���Eb���(5DaIf;��}opn<D~����D��F�`���s��s.�*M�ܺ�BG_�
aۺBx*nP��ǰ�4kv!z��u@,�(k� 9�/���)�#_�..m����2;w�;�L�uT�?�VL%�<O� �jv�"�J���r�kS��-��X,��a��s��%���s�Gnl�f�]�,�K	R���#� Y��bV#8������ќM�"�L�C)�YX��c��lT[�/(~0�L-�4�96�VP��-Ud�7Rf�9d`��߽@	��+z�_?:�;Mq�� f5DO��$�=b�v��ſ�P��KVA7F�����~��T���2N��~�0PE�F�O�췢6L����<�nw�Vr�S�&W�ϑ���^Pa�Ą�sR�������jf���j�<�p��(�'�4�Q��zZ�c�̿X��F��7[q�U�~@t����w����$r���=�S�=`�. �2���i;W�7N�wD]q�����Tz0
����O�0S6U�KQ��j�KjQ �LP�17�|p#��L�ɏ�@=�����?Pѹ^�� ��b�޻/8�0<uS:E�;Nw%�.�u ��椝�w��3���MI�X��h�L��t�)���i1s]m����F �C��oq�F�9�qh}J&�s`�-P�N��Yw��'��YOM��y�/F��� ?n�KŨ��=[����*-�?M3�+^Jb��$�i�����M��u;��~xJ�`'�o����������a�3���2��R?���������#6'1�"<|�:�%F�`���	�h	Z;VmxC���#rbR��O���4O�3@́֜f)�?O�vm%��Ew�#�����ϑlQ��9�J�&^n�_~����G��$�%���R�N=����H�6.M�Vt�������|������}�#�4%������XC���@���P�뢒�AMӏ�2��<݋sv�⡬�:�f���%߬�� ��*��b�r�N8���7/{��I�8W��r"�3�xܱ���ίw.wH�|��G�m:f�LH1���F�.��]�3�0:�!>ÏZ�ʽ��J*�~8�=�ο�rB�G�}�1��%��uci�v$z���|���ypq$q-t��V�O�րB�v�9���Y�:��>�VyJ�W173[�ĆG�g��YԺ��S�a�
=f�ik�M^��'�\f,�ԟd�Z��	5=ͱ/I���b��8�|:�.(���(��v�E����\��XҶ��ҝA���Q�d�j�D�:2�x�Ǉ/�ƻ���e@�L\�t'�=R��eN?��LX��͉l_f��_��]+δ\��W�Ye�Y�C�-(,4��7-�2u��5Fż��}�%w	e~���# Nt��6.�������NS��wM��:4=K�z�2C�5�Q�_�4��>hl��\\�M� |�2�����U���㙺 	��3�qC����j+Wz��W��F�B�@k�qCC��|��?zX��y�_<l��8X+X���u;���!	��|/�~�ƶmۈ��[C�����)[�ϊ�z���̹��8���KՊ�@5��Q[^8
�\baVH���XQ�a`X��PE�����t��ZrD߇W7̣�ˁ����&2� ��������sZ��.���v����TaHQӈ���,��$�J �zМ�P �ߢ�[�}o�io߾dh������y�����ϰk����N=��a�29J���*�ts l8�(���q����!0;��E�ʁ�ؙʡ����	�I����b���â�~���/E����ViY~
ls��r+�q�ن��  AT��u�"g{m�&�L�?C���H�{��6���j��:���FtB�ٙ��D�|#�fw )�Qmz��8��afp�0&�Gʫ�h�	��ʋ��)�JY��Ճ�΋����[���k���i�����֤�*Fk@�gmA��{0?
�z�� y���K׈���0Ú��68�v���61�C�c~��c*�'�n��y�FK�ݼu+�2��e(��u��3F�nTcO{(P�{��G7gh_��Ϟ�p�O�8z�Dό�	홹]�q��b+#�aڻ�(���k�_
���R*��.���G��~�〴�(��܈����^G(S�n��M%�젩i��˗/��}O���-t_�vm�SO1�>3�عx�"�?�o�4t���u�D�Ak9�KpT46���,�UY��[dj�����kY�mО���TS:s� �Z?9��oP�1r�5���;�ewLw	<l�� ��6�(�x��L�����$aإp�So^N��5Pw��7�Q�������:bL?���D���vgݻw�����o������)� �5#�/�F��|,͍��2
�~�c��d�;�/�w��0E>'Y*͡�i�d��? �k�N�
'���+dj�9�ɽ§��w��a:�@X�j�+U׵��z�
Lz|Y�B^�'4l�eS��M9�l @�@��וz���^l����>�Q��o��B�`w�b���b��2�[2zf���^�L&�\�{����[��d�����aܳ��/��>���쵈�5�S���d_�:�鄧��;:Db�^K���])C� �~_;\���k~
��X��BOZ)���ĜB�6��whWMۖs73�|�Z[�^ ��lfH�L���;��H���tJ�gV~��dV<���~��0�%>�WL���kV��FIw���FO�+�\4��M�{gMF#��cfӑ�S�2���7�^ݺ�@�����"2�Q�'��ǆ[q~�}Ip.�'!��\�<�n
�W(9]1n����&�z#��PB��y_� w����Y�^\S{��}��B��u���=	�̜�{e�cP?��z�k]��B��g3���2�5I��L�\�w
��I�m��|b�Se�Sm�~���O.lB&4ۼ3�sW��B)؂~y}�^�S&�b�΂�RW�;��|�ra]��i��r�k@�OQ`���"�;�I��&�4H���ʔ�_?�]{�L�1gϞ=S��i�����5�)�E��c&��dcgɵư���84J��N���f���Z�+A!��n�|˼#��n��O�<��}TS���YY1�g�.�V� 1� ���N}��D��5J:8�;� F�b,�-**JW}�N�OjQ�]�p#���x3���j$�A�ry��L�������ٗ%�- �f����F�c?+���M���n��:�U�L�	�B,��fJ	Uڌ\/	2����u��bX<�^<��8$�I�:��n�n<n��%֏C�:a��	�O}��%��G.{4zrL����C(��>_x�+��\�%��I���;n|�{\���~v '�Pz��{��޺�۸؊3=����8w�.'XrQ��p&<Յ%W�o/�c<G̢�_5ǂG���+�yV<��C'��[�f��{������h����*U���o�F��`���ͼ򷙼D,V�ň��d9���^�B
͝ȼ&�_�w��	�\/�F,�	�g-�0��}�di #��>�WRW�3��irdw�H��#+�H��/��N܀��R ��b��(�VG�V	I�y�z�{l��K�G�5d�ʟ�_�3��Y����Co�c�zz��o��Qڈ1$x��u#�C�>����t�4�5_�������526!�=HƯY@k�6����';��)�b�,L�il�VwZE��[O�3��g�7v=}�tkϧI
�<n����~G���΀/@[���d��1�ӈ�|�.S�9bs�`qp��O��Z?H��\/���I+ŀ��>��FI�3� ���`���1ڒ�z���`�.ؠR�UC�й��.�+�@�'����	�>��.v#ԸSV�<�q� ���S����uz��X�{��v]O��f�Z���=����%���*��Щ������������e���}��X�O���f \��+U�:WNw�������в��v7�im1��r�CAq���d�ۘ<ώ<{2Ԩ!�w�ͅe��f��ؤ��/�d�K,y��9u�=��hl��G�t�W��|��fϝ��`�k�`�0��A�l=�+v�}�6����'�JmJ��+U��I�q5	r��E΋�z4�*\[w�'}'��m�o��U;.���:i��$����{��'��w@%��q�{1�s�oL,�Q��s~#�s=�� ����}et�Z�Zw��J�?eKa�2���pGlC�}!Y��$��t!�G���a	�))�������\��~~S�7SRxv��wPj��]�V�{/��`�-�o]����H䅶�]	���DZ�f�;E�h�����:>�&����8: �I�c�%��0��0:%C�7��c��Ka�Z�0qY�/y�8b5Q���j~��Z�h'��!7�%��M,�2�簈��������S�]�ČRC"�6NHt�:�Gzr��y���rA���
�C�A�ȈD���,4u�����e��w[�Cw�م	,��}�b�����`rr2S:�����@�;Wp��#r�l��O3Ж�cF��ݔ�x �����֔V�0/cv
뉬[�=K�ӟ��rҨ)�nXM1]kt�燌Mٱ�P|/������j8p��&茺�D�w���6�(�4�9 �f�#�k5��.
���^����j͈8�f�����B��K�̓�=�v�\z�R+���I���v�7��a��-$�^S�b�*}����>�&�E׳2��%�62ed3�0�i�51��i�Ob]�c}?�<���䥘�>���}f�	�}^n�B�n��o@'H��Dq.�������`x^T��@�?���yϦ�E�vj��q/�܋W��Bb=� ��FǞ;�r/��gg
�'��.~I����k?P��LdVN�eB��`��6�R���K�mb�f.	�h_p<ΜȌ�I�p�eJbZ��$���Pkf�0P�K�"�l��n>xY����^��Vi��l���6.f|��Uf�]遗���n����/��͋���0���r���Ϋ�1,�d��{�5�����+��[H�����		)'��/��a����r+C����ġv�"�������}�0���-�)�lKfhU�� ���r�j����	�]�W#!CD��a��ń�l��D*�J�=T������=&P������U��ow��H!�)O��Q�Xm���|o��� $VQ��ޠ��b�Z����/:u�C�!���[�4��^��	��:�mE���7�H=��/���E}3�J.3���;�Y"�^�R(��7����zP����j9G�&'�r�
.5�~��
�������{ٲ1�L'��[ųQ�V0��a�(�0썝�F�ڇ8pT=�/zC�"7�N[���Q��755]���
��{�]�F�ͻbK��۱�0�
���NK%�����IO}mo$��.���R�k���|��LO�����5l�0Z*
����wPN���%n�����g�=e�tP�;�οv��mz�j>�a��bx���W��®�@h��o�&�۱k��SX0��b0Ă�L������������e�5>�7m���d�ơ���>�34Z�Ʉ�r�fҿ��f!&|�Գ�~NNNW �N���0r���<l_����'���b���!Z"�����b#@l6C�OF\�*	�#�c��P���٣��p��K�M�a����]���]�1&6�X��)�-�v�X�6��r��g�]���Q�|:v�>c�'�}5���(w[��-CB�@"�̖[� J��D��j�%�6�kn���a<�/v~�r�ޚ����U8ه� 2I�.Ҿ}�����m �9�b�D<�:/k��/�EwL�!P�|+���A�sJ`)�� �te��);t�frՔ{���xjZ���shttt8�r��xr�v\g����<^�ܰAv�> ��n���7� ��o
��H��mL�ڶ��N�30�����aml�3���u�]��(H���&ƀfkx#���.�Ef����i �Bw�@�?R& �;6�V�<�����%x�����<�M�L���1��w��;�JXn�uA���g���K��Oa;�,��~%��#V͆k	�h��}�\�c:�j`XgJ��D��_�tu����%ڋ+2��ȉ���*�Z@>��Ø��2�h-���1�g 5��_'�jFt����̣	j�<�w�չ��T[�_>����:`��w�~�u����@⯵�;B���FW�8dn����1U���R�/��En���
m*�w]�r���հOnq���?r
����x]���Sߝ���yݬ�nS}j�r\�J�͙��;�C�Y��e$��!��8�$O yݼ	L�F�;����x�ꗒ��z���~��*������+7{x��s�0�?�+���b�<ɭ���2�=T`�F���C?YB��5�¡=�V���Z3���E��׈���&��҇]�j��z���0��R�
YulX�J��!0�H�z��i�O�g������{*m�ּ�M@˟���bʟ|�W�cV`.V|1gOݒ�%�(����3�B�7�U$�C��w����5�Pi�u��
��B;�5i����M�L]ҙ���������������u�@�s���ߤ�@1f�y�����5~�:�'}�탕��F2�KS2?5�$�oO����9C1e���̎�L�����f���O�;��g>3��jD���*:$HQ�yp�;	�IK���5VJ� ��{[��r��_P��d�͘�:���'��d___�4����19(�C�Ńhʩ	�^P1�>/��P���;$y?����1��yq=QԊ�[��=;�lb]��������N��%(��LA�E��Q�J�c�}�i�\+�3��Ä�z��
G�����au�O͒Rl��q[x9�6u��ӽܡ2�Y��]��OR��-]B�5�\��X��7jrU�8<2�hz�BGqv�+Є�{�k�z�\�2��5�ĲC��Y�:g3Me��v��2�,���Ĺ����Kw����H�var�x�!_�7־�Q;^ߏ�-z=�k�L���D�**U�����VZe��<z}d���xzK������cv���MgY���d���\�J�}|N�����~��}w�cφB0co1�	�Y����2cv�Y���K�M��tp������j���I*�n�!!!�D��kmGH�%<�E5�f*���m@���:l��zs{�y����K��0�ѷ	Ԃ�('�'|�+)<����g��Oz��5��e�j嵅�k�2U��� �_Ǳ*v
����^#f��H����hN��PC�#ƍȤ�X���@��vIp�$��u��ܧy]9		�"s�ZO,&7�RM&B��<w�OM�e�L���m��-C��4,��1��&\�k��]7$�g|T5~y���N�n�8妀�����Ж8��o~�dovv�­��㴋�K;p4���n[^F��%�:�=��H���yM�8����YZ�ڊ�˗�߲P���yyO*+%��)�Js�%��]��6_o�|����MOn��L�����t�ȁ�EQ�x��{�c���E'��'IJ����-�ٍc���5T!�=I�:�5��}�"E�밼�����~���u'�I���C8Qjvy%'�M�5�}%��|�z(�?ȫ1��p�mb��$�}D�$o���]�����Ę�q,�m*�Fŉ
���cIj9��s�j��Ir*��֛$�b���0!O�Q���G"Ӄk�6�4���<Q:�3�$`&;�I�4��7�ԥ<��#������)@��?yr;QZ^�oT�1���T�CY	9�,�"4q���Q�ר��SQ��??���*'�p��;�	b���SQ�}
�V���{�n����Z�[@�^���֋�,*:��=���/\��.�f=IM�J��{�>sÆ�qP��E^�J�[8���#���O#������D�Yq�p��~��q�6I8���ar!�SǪ�'qo�x�l&a��0d�xJ]��cy�jl,9�HA⺈dyW��r�ti`R�h7����������wČi�e�t�f�&�t@ZN��k�4�Xہ�1�H݁���X.�\u�RÚ��]�ݛ�bs�&��ƀ}�*��͏)QIޫ���i�Y
��O����V����@�&�A��9���4�c]d	߈M�$8���fh´D�-�5n��hK"�d0����>\O��m��Xl툺,�2]I�/�7���IB�%B=�z �$�p��0R�NI�+Կ��bh�i�ǇIR�h	���Ƚ�L5�ɫ"��Z��|^kf(�l���	������8��.ryq�/2��?���p�&�w�9� �R��`����.��*{��Y5�/XM�_��C�*��$����$�覠���  x���#f?YiI�Tkex��;�,�b����zJ�)�>�M��I�=�^c�C�hb#�ʂm"-1"k���G��ʊȫ��q��'~u.����ƍ7����]A�զ !$>�J�l����0�t��O�����~���Y��r�@>���Rjm����G�~mmm]-	o1l��E���."W���8c�MC�p�ed�w�o&6i�$O���o8<�m�!V�m��w���Ν��/$�?	NB�Zci�.ߣ�Y�r��J)QH�8Uň�#�A�5��|�z( %=�����r��N\mxKU,�y�=���v8I���V��R�'Rq�x��|�؈kp���4N׎�m��}#"�S%%<0���߲��Q������8��\!����h�V��m�6�#ݦI!~WK�WD���Mݴ��*��ȳHOs�$ʛ�3(���d�K�?L���Y����H؏�d%kV���>Í��>���|��7�I�B��űv���B6~��|[��q`&�*��6ܼu���\�	�9���<K)!�=�gy�v�&{�3g~D�撤t�q�7 ��G���~�&��NR� �%��.�b�A�&��ִ�m��`���C�Y&��:Aʈh���n{3`a fՖ���4rn����'&�>�i�"dnǥ:�;��v�Kޝ�'O>1P������{i�S����d��[�閍9���������̝�+T_Ϩ(װ�&*=-��=4"�!�T�2�:�T��$�aN�����٢G`#����<$��L�.��G�lB��-�]�T���*	��[;��!��W
��2:�pO��HC��!��p|�K�7NVEJi�����u�W��B?��FZ�D��L/���Px&D"Eo)vq3j@,7RU&�>�ΫKsa�yi��m���2?�a�Y�۞n�/�ޡ���f�ǩS�΄=w''']�^�;h!)��h�MF���_<~xc�u��ŻFQ�?~�tɑ�4�\Z�s�j8�.i��(�]��b�j1��*�Ӗ�-�b˦�>˛�Ns(�$��˽;�?C�5�R����Pd�(�겟�͗?�������o�$Y3׍���~g""=S�*�y@]z�c���Iv'X�onnn�Zk����dz��545�%$~��h��!�t��w&�<��u�Z�C����r�����]i��8��� �|���U���O�v,	)ֵ�]Mv����W�\A����ݮ��<�U5 �!�N�c�Iᶢ2��'��	�c�y,��wi��oh�N��#H��Y�� ��V�oDF����V���Z�y�Yic�����V9��D�ѣ��
v?���;�x}^���J>��6�|	���QU"���Y��?ۡ�Q��S���\���G�m? s*=��d)�;�w"��ݢ�Dcp�Ν�tL�3����T���#v����D�0���0o�-� G�����'~�V���x�('2[�qFF��pcC8p<+YW�e�];�|z�����b�赞�

��؁99&؄�܀���/���bAK̐5���[5��e2H�R�Ϟ�)44t�ə�>��k�= kk-ށ@�aR�e�h;v��g۪�o>|�P+�;X!����	�u-H�濔L+�*QhN}� �OL�c���X�ہ�T��{'�!��
Ę�a�0�#.��sU��:����2D"q2�.#+������*]�o��/B+#�dx<��g��OU��xO=�YN͌�E����	��

A���5�F��S�Q��������,*�����ۀD�>G��L�Sw�J?'yL��|\\\ijH,�A�&���"�~���v=�
��X^��b���O�\2���*��@���8JLL9#?J-ph��՘y	m���[մ�ZS��e����L YH|��cPx�!;Ā5��`̈́����>Fm~���\F��G7�� .j� ֓S��$!��� �����}��6�_5�EOe�`�pV��,�ʖ���i֘ �i�JI�9::�/*���֭���6�DG���w�h�� g�u�	Y��x���Ԑ�B~b�XzN|ej�Jr��{[GL��cW؋$5��cv�i��zN(LnI�sL��@��hP� d�WC�|���@�)��PU�[tOxS��,//�h��օ[�� 㝀,�_�u���.�c^�^π���J, �\�����+=}}��PUU7@����{�V�W�
��lSz��|�x��U7H��Ջ#����tedd�#h��(���Pl(���b ������R.�Ҩ �gQ:J@~�
�q���5+��R�zzּ��`T�?��Qw6�(�?=Kw�LN�`@�(۫I����Y�D�l�����BUj�/B@b#����u��s���UTz�.���S���T��>��}ܭ�����R�n`���Χ;�{�]|_J��8P��NV��������s�� ?��th7[�֜}��*P��?S����'�o�����ۋ����Q̪%�Z�J���d��'���0��֣��¨�{�|�pVN��= 3���p%p�,��?�G�c��~���y����������{  ��������Hi����b��X�@E�p�r�wՁ4O����������A����>y�ys|ǡ�WQX����� �Z�bd JK��B����kV��o�w�n�\���u-{��˸k%Ф::bڲ����_=G�����B3w_��+@�;#nݺ�`������y~��[���C�r�a��$�`���~mo5����C�� rZoo�9K����c��z�:r?77�Nk,�6X������W�Ԕ��G����$om��+A��y	�q�8�E ��a[.c��}�!�>H����D0�u��볏�vQ�0��ͯ���h�g�B�Ɠ�0�����v� ��SK�L�Y�G#�w���#diJ_��2��� P�`=V���Z7��E�oL�*!5A�s��X�/\k�G,i�K�R������	D�i4��Pz^eô,UI�U����@(E��a��)�[)���O� a�`-�B�>�-�T�B~R4��"y9	�f�)���i�	�O-9��W_9A��k-MM��8�Є���%�P�2 �ҽ�u�z��o3��VA9��1U [O]��f��E��ٛ�@��F4G;� U�yz����DϐG=�p��s�As�u�Z��*y@�21q�4�,���~>[:,A�jڥ����7/Zo�읉�73c�����k����E {r�$�h�VCړ��I�U�V�vj�kf`U�F�	�x��ъT�c�lA�1�n�3�o߾�I\Ɲ|?	`rz�8绮X�,��h"V�Ov�Ծ�-� �a���e�agg��Pe�֫t���u��9?�$���}�NG���Y@7
8��~��d���u=O�w������Oh��)v��I�?@�;W={13VG/q�*E����W('M>ɡ=@������g���u�"��;�5ѝ=P�����70f�����Ѫ���)�j�Wfǭ��/��I��-j-2Lu�L0��]�* ���	ľ�Ӄ�݀%ש�m�%(hh�*+��H7��k�ĭ�1�4/[V�!纈 ���6vv���X�?�a�Q��n�$�l@�t�իW)�5�;���n�-�!cO�� ����%	M�NB��z��m)��R��C�.���!��D��{)A�g£J� k?�������])�)���Ǖl�g��
���ů�aD�
2U��i���6�b��߮��҈�H�]�R��8Vڡ̬,���.0���7T�t���N҉��Df�H�����r����B�'�����';>������ۈ���xfcqq4�I���,P陃Ue�P`��%�cJP۵�%!R�O�4��H��ȀsF�t�Ò$k����K��~?��\�w���\%;:�C��}����2T�3��*v񈼭h9?�v8�k���sp}���~�uua;6zz�$h����M�%�{$N�DO��R�Lq��Z�v���i6S?B�lY{~��ǜ�ˏ]�x���WS��!�?��c ���G�0�1G�S_���p]�)�8V��O@�lml�� �\/�u(�~۰��o���
M���͸�Z���ΚY��YY
�������7ե����}����?���g�����|�F~*Oc�Z￀�.�,P�����EYr)VB��moVI;fm4�j��g���@��q����s_��'�˷�⦥�.0+.Z��}q ���F�(��2m�S�	���̈\ǃ���2��P�4/�;J]��A�#N5��fv��yg��?�Y+�(5��v�o>���@��m��x��-,�R�'�������{�� �DjZ۹ҫ-Ye2�dߏ�gdK����="d�x��I�u�,϶@����߲f9�_�ˡݽR��e��T��Kx"`��T��g>]����{�A�O�UkhxO�g�KOj��[f*&4M���4����NX!�QPX�<��PL)5�S�OjJ�y ��HNIq�f�#�EE� ����J�����6��r��y�왯o	U6�V�4,�z/�t@O!�P�0�PP�� ��=��F50�,�ݨm�\�%����B�	jCnQ��S;7nQ�>���|��������Pf�o����I�]��ѕi�(z��'f��i|���	�A�w�Ø��&����%b��^ ���j�ZBh��!��,��

@υ#��-�E��^�(�(CrRg��"�&�A�~���Ю���O�g�qu��m
 1l�E#o~D#)�Z&�{?�h��af�� c���r\�"� �7IVA�$+-�Ut �xy�^G���C�`�o�k���eW"�1?uP����w�T����ű�� ����|�f���*CD��]�a�/7��;�h��T@]*�;o|�o��s������#������k(}dI��`��052���c�%F�I(�ۓ�Q�k�$`�ÿdkV�6��m&$~�*dl�+wD�W�+�k�4U�������/. l><}�7�����Dy�#������)�й~��\�vє���"��h���pav���"�� ��k��^G @�`���~([3�<6����9�뮃��S9����Y��O�7B��t1U��N@��5�k�B�<(�`'  ���X�W'�]m=*��R�^�X)�f��5"��  �4��G1��ф���z��oP4��QZ��By'�Ҭr�l50�X�׀Ð����ue=q�"c�Ƃ����/�o���-WT����Iȟ?UiD�j�9�2�
J�r�@���4��������"��P�'ĮO���~��a��Q�
�1!����0���zP8h��(�a~�ڠ���=��D�O���\m���h+��.$��|��b�.v���В�SG6q���D��+��j�Y�����G���e� J�n�?�̆k^�z��)�j"�	�{�\��#U�5vQ��K�_ׯ��)��0O�Mg�Me�0�`�)7��d��{n�D�3�'aK@o�q�=*���̊Љ�0�b�!0��vG���w8D�����k�������&�^c�o:G����ˣy�90��Y���x�-�����	��=���̭��2�Z���*��[�5�/A�T�_o�=����^ ���O�G�W<sZ��o$����ǯ5U3!k�_4[��:9�(>�?ȍ攫^
��O����p�F ���fh�+��������W���^����k~��Ly$�n�\s` �@�=0��s��,�GGyG�)��mC�* �V�"�qB�Z��m���w��a1q0A�:�˨�uؖ��3�4 �/hU������ �r����8-��l�J!22^�4(Y�d+�M�^�SVHB�5*+��{UV��[F�����_�����r]]�㹟�����>���s�l⋞;\c,�ӛ}d���9��B�г�+f˃�r$�X���lV�~�����Q?YQ,�cҰ;ТQ*���R�Bv��/�yyy�'Q��0�m��O��.� �ߠ�j[�����~����1��T�*B�ё���Rav+	27���O���0�z�Y5S�}�1�L;^�3ˆ�)�B� w;���QU\�[Ā�\7��_��2����ō�T�O%� ��#��o3��ބ��ɾ���_� ��y�8�����a����DTV$E�Ë������О�I���nc������9]���F��%���9y����&��f�+�av{��������c̫�vW��t	9�E��'�~<�u�vt��x�<0D�����?�N���9�Q{)^�~��P|S���]>`$�I�ɹ�B��VQo���	���{1�/�k��3:::�/���}�����I l����j^-��`�4128�˟���`�k���@��bڹt]�O�����ׯ_�S�V5���	�CCC�	u;4QUIde��������d���zy
���p8�d�Y8El��
t��leuu3�}	���&obb"%%U\T$6]|�/**j��ډ2J����]W���~�)m�{K����p�J���Vښ��W�J�2w5���Z��Bwإ.Mܖ�i��O
��������VW�l���v�I�17][�n@F�2++��H<���N~d�]��K���c�q&>������:�iu����}��FI���eJ(��&U�k	wn�dV���x�1��n�U9%��T���c�(p/%Gd�(���	;�����wmy��e�L탛�h5��Tt^�re�⩍Ӗ7Y-��˖�l:�^���jְ�`ee%��2	�U]�y"��5{��u��J��ˑ�\���
循�*�P@J�ǥJ$b7!�?���?u>N���2<���L��sG�:�`ĺ�����E����p��)t�,e�X�H�2Z�R�T��|Te��TG����ġ��n���O��4�@a��C��P�Q�!��3�C1m�JDSS�H��*a�FZЫ��g�K�[s��4�F�RŴ勺��7�z���/�G��kH222z�4������kLyQ��(]�گ?-��KY��(���yTq���P��4o}���
�W���KPWv{�wKB9��3<�֩��|W
!q������@��}SS��
���!�f���69g�w�MHꡃ�����-,D������>ׄj6�����.�rN�y�Ǥm�>�:αa���go:a^T��A2����}�D�c
�q�����1q����C��)�Й��r%w�x�>��&�
� ykuyzE7m�@��=T��@�op����Ẩ��������9Q�}q
����l8g�t��o��$��l�����Ə�\3�&r'���ofȝ[Ӂ����𗖕���g%��,�ro�����T����'��JK�tʶ��b/�TPP`������P�p�x��d��hB��V��-;�*��uĸ���F>[�ƍ�s��z����J�?���r��>f�������7�A�nB��]����3P�������m~�
�K�ӗެ��`g�����oE�-�]���>o�\�7@Q���޹��41z���YT�Pq[|�+���w�Q˳1=Q����D���X����J\JN���W�ޮ|��,gD�?��(�ɲ��Nc�zո*dqn��X�N�h����ڧ!�Q��w����CօG??=@��S��%��>���-C�%Y��9Q�+|}L�Vm�x�8&��(la��D���q>�}��5��FȖ	��GM��}%�5����b���;����i=@��M\��Tmc#��t��ř4�^^����"U� pa���k{컬fq�&Ϋ�+=��8RL7+,�IF�{466R10�LLL4�%��(�L~���rW�4��0�+�nß��c�]��g�
��sW;,B��E�iM�}�:M��
h��}0����^�:��Ǐ�UVS{θ�T��)��w�������?J]��̉����e�D���l��ᆠ����iJJ�m�~��b�U͔��x��տ �N1^
�̲���`y�*ȡ*<���I�pZ؈���r/�����j;8���mA�ϕ���o����*���A�-�����qw��(Agno���x��VE���O����(��R1�u�gƣ���!�F�X�t���V� "�g*8ʼi�vNL'v� 5V˱����x��x7hG�x������@�eϠϹjjo_�/v���|�tj�:�����C�E1�`�^���(\7�}BJ�p�XS�������������o�/��0�2���������s555|���&f��V6pbҘ�w�v� ��@�vo	������?{�l+����E����ܐ;�'E0�y�/���{��#C�����7x�;���+�
(�H(�lg�%Х�S��u2
�d�����a�1.L)�w��j�%�U��M+q맷���WVVD�#�ܻ��|8(����A� ��N/���+R ��w�ې�n�&^��ݦϛoa~a���Ԇґtt�=<<�&&P�|����[ $ 2�^V��Q�at>�Q��N<H,�G��sssrr����/�;{�w��|��5vwo8O�h"���gA��~ӈ��^@e�`Q �/S/��UN�s��%�39 �nBn��J���;��:��)���3ww3C����8�9T͸��K��M�:�Z�ߚ��`t�]i�Hd`F-��]�cQWW7]k������x�J�����&Hy\$�=C�4����@��;T���ۑm�\P��`�kbW���7�7�4�x�.2��"	ג�=���S�����H鞞�����n��L��5�U`�a���d��m�S��o3�5��S��-#?�~�
�500��� (;�D�UM�/utv��O�� �FA��s뼽�t�ҡ�C�ng`` �Ծv�����M����Ɔ/���$)���O��]��k��nr��3��Ҋ��֒�Q��bW�p��5Y�^Y$��T�p�
y�n���;w�ܷ� �%�e��xҞl���:���E2F�w��qt����{�yB+	�ʊw[��/�?��,�0f�|E�3%�#� P�gϞ����E��1�3���|�ŉ�աx5������@�>���Z�#����u���wܤp�*ou"7�{�M��4���M�AJ��������Oʄ�л��#$��\y
-�z�����������W���վ����	��,���_
��I��ʁۥB���셬�^R��ɐ������Qo��8���1�nX�؍щ��͛�?�K�����:��W�Ǆ���nN����b6y%�5889����[�w�Đ�>zmbd4^}��Y
T�/_8ED� (N�%$$�#=}�4�r4pt,�ﴶ$�I29��n3�V%a[�E\��&���V��>Q�X�ӽ��`ue4a�;T�g���C� �_`�`�(j�Ns�Z��v$��&rbk���ٌ����' ,,-K��"'M�~+����{'����jd��ݏj�Y6�?�l���[��x"oh-���Aac��I  3��[0���C(�}�����|轠�`�S�Ay����2e�<~�]��{��FGW�RV!'�A�����!;�=�%�jW:k��8\ы�Y�񣚔@�@t�c���+�"�&b#�v9��pjh��f�o��^�w�$��������|cWX�5�Hl��9.�&���v����E�8߬+W���e��D�B�t�����!��3����}�gΏ�#��O�s��j$ߖ��o�D�-�\�	���ZX_OJM=|���w<Ӹ���o�=((�7XK��0��Jo��@�U8��P�;�#��ZD�u\�?��>�{l��Ī*^��6hN,���GM�+immMX�����7H(�HK�O������2������ �c/o����v{��������.M�Ak��5�xM����,���[�i��ɫ�iQhPVn�E�$Pr�M]�(p��p\�h��QPQ�L�6�iRS{��T�+))�a���8Y$�k,�\�ZK�g������;�*�Ht�qT��W7G���U�G��0�3E��^+P�����ؽ.d�YYT���(��w�MQ�F���*���������{���A9G�jNh(����zH���q��@�'�$�6�+��/v�" P�Zѕ��
�}�ɯ��<4�}����*��E�,ⴚv@�JJ� 
G��T�B���'�AA}3���G�s�E?i�uˊ,?pX��E:]�t8_t
�n�3�*��@Џ�͋&)l�V(���
12�"{�H]8��)�76�J��"!l��U4Bw8�y�t�#;�|PfGZ��-�z���E��"�DD6b(����A�8&�re4nn�)cV�@�Iw��H\L�pL���*�qd	H$��sS��6>�d�e"�	�)�e���!���P����8�@��
ٽh��~���P����%I����*��RQ�����E��Ӽ�Ꮤ&O���J�� �!:�Ō�t���%%�A0���l�G����ܔ��`�#,�et[����Kɓ��D������n��I$" Q��Ĩ蚛s;M{i��Y(�76��҂�C;�nP���Z��J9[�g�ys��$�&x�ʑ��E�C��gݗ�A=Z���7�)��co����8���84}���aI[�,��/�W-<V��^��n�y�51��΢���qT�/*�q�p�>e��ԕi�)4]|��&�^d}��b'V�f�-_VVW�PNM�fCk����n�)))�E�>����{���D��<y>�{J�o��8L��������Z�a��d������Y��#�[a�{�w�WƖ��^�D=��dٽ���g�pa}cjj�_]}�&֘746��Lc7N�sv����$����5�܅���W[O��R�T�KS?�+���&;on�;,=�^Yi�U��o��		��/��-�.W$�IQi��*�Rhu,U=J~�:�q�[CY�*]BSSs�c����ӭsK.�����V���7@�A=��rC2�"�C�j�А.�����c���Uv���*�!]�Ųq�iѫke�?A��[&����������θ�*�)��E�$����@���*�����Բ�΀c��u��$�i�D�Бz�jΊof���C�8��ބ&ˤ�x�Y�gXXX� �A2_���`��`�k�~����겎5dP�ۺX����w� w �Q}z3͕�&��z��2(\ˁ����o�$A�K8;;��a���N>�Q<?ڌ�F�ҿ81! `i�7���q#`+o�����.���'�Ք|�Z/ҸT���z˨H�_TTT �_�:YȈ� Y�񶎎�qqqw55}��;��:<�?��F��xd��c���a�N�-���5:hk3���}��sQkmm��\D�{�=�Up6�[������Q*0O��Yr-���KI �����g.����|�!�vzF::̀��p����Dc`�&7��z�L��@~�ZKq�� �������Z&� ������o@�K%��zO��v�D5v�(����g����ϓ��"�jI&V�k>XEM��>
��ؘ!T3-���B����o���`A��=D~-� ٙ`� ��s�� ����^�`QI���h៬�A�B2@\z}q#���At�8'��v[��I���w��J�f��,Lv3:::��0v6���x������E���6���$b��(р��ST�̈́�I����;�P]966Vܙk����P�.B+�u�Q�y�)�\���ML116.���s�x�8��6K��l%__%_�s��,iDԷ3)YY�H9w��]_?�Yo���W�Lj���)4�Q��%hC3��6.�H��b�� �M=�� �z�9As��+�m��jl��@nף�H���r38��6w,��G+��>��&5$��t���=n�_:Θ	P��F��>
�x�΋?��4解�a�"��螁ktt�[�:��X7T[>􂔨��v�JH�e�{�ZP2��V��*C�c��i�хJf�E8 J�M&����ʥ�/�} Pk�����ZZZ'��V�Gwm.h��%ݔ�i��@����P�������u��Q(�4o�#���Crj�?�4!����R�[����N�"�� �v�B�Eڊ�L��l�9(��Pȣ���\\����&0h<,!�r�l
�MT��8�7���ɀ��ז��W�ve\`W��4�{z}�z///�)��Ɖ!��h�A�"�9�epx�/�`�ʊ��Qa=@՟��}�~[�\�E�� !턷�W]N�`"tyk\h
ncf٘u��2����ũCp2��`�C$c�R�jp��8�%:��t��o	�a�]#�����.��������h���{hӾ�����xS10TU�?�Zp��Y�c��Y�r�X(f�[oq&(����x/AL+q���}��࡙��J��?,���M� LH	`r"	
R�č��5vo�v�ҙ34��08E������i�pь��_4.y���W�����1E>�*�Ϗ��OG0UVU�zqPm=MĶ����:	#4]__�мB.ٗ�l����0RH�Dq}kK� �! ��e�Ƽ-�����7tn2Q㍨�H�t!+��S(�FH��K�� a�U˷ۡ��{�dS�������a�� �����C�K({|ᆝZ�Я�$�ddd$�Ő���@�+q24>0�����|Ң�vU�����1-e*�F�{���A���&��B�8C�{Od��y�6�A�$k�ՕN� �w�����<6qS�=;�5�p�����������#�T
�ךlik�w�������#��d3���e������0b̾��@ƠG	=t�٧O���ǥq�S�	������� ��*��:r�9��kME�<8�
��	 p'(�!(nh�gv8u��~����V^��&B��^�s�NG��~�kJB���]�r����G��i�j&��;���w����L�����_r�(䏉���j�!�P텄j�¸qqK�O��6��g�F=��������넥]A0�`4��]:�t�x��IgǺA���z�����o�{�#�/pp�!$F��Y:%���V��dcamSu�� � Ը3��C"N3ҥ�����J�7G_A��U,�W�p�Ҁ�� h�t�G��j�M 2(!4V�{�=U�z%8Eꌻ����6�
k*�i���̸��ͣH�C�HZ�&g��K_b���l�TUU5]]'<����ߗg�
�����g�3e��=|SX�t.o:��32(�f��nQ=7T����		%��f�E�6���iP�}NK��yP�W���3�m��r�"h(���Ω�O������?A�CT�,?1\7@�q�	c1(W0x���cʢ���b���áw� "��٥Y��\��V�C(m� ����\�=zb��q��Q�/��ǃ�Dϳ���r�|qC�A��<�5�,�	x����?~t�E~l�GJ{�1���2��lmQ�r{��q�K
f&���@#֓];�最R<]Ũ2�oCn`H��yl�N<���E>V�V���ٞi#C�u�z��j/abbf�=Q-�0������lcG���6P0T����l]II�Ɔ��iW�	?����c��W�[A�11
:��=h~A@ݗഠ���]�yn���_���6����'̡b"x72�G8I�y��iq48]�����4:z�o���;�Z::�v��/,�]:��T�����ι��a���&m�3���J����9��.Bq�t@���|e�W�J���}"��<#>!6�;�AGb�1 *�ˑPgF��@y�:xSD�
��-yQ��`8��/#��h��lg�/o�Q`K��"�r����֮.(R�x:1�Ah 9Z���q>Q�B�m��> ]q��t�v<�������t���ߒ��M?Y����� V�����Bd�\Aq�GNJZ:�
q�!e�	Cؗ� �)(���^dm��z�s9}�yb�|��볝�vTN�w8�|�����'�R��d?�v��yL��(;�h0������
�1�r;Q�VG��V5���e�����`�F�2@6�����#uޔ��#P�28l �L&�\�v�]6GX7���:+?	�9�!>��I������QU`u�Hcvv6��{���Qȃ�Wv�3U�;��%���颭%������+�����UWG��	�6�o�����)�d/Zлv�?C�=��;bw����������X?uxS���+�|�SC�"�R��^\II	hN���{@�Q|a�؅A�I�����j�F������L=�S����}���L���1)���jW�.O�Hc|rZ�+lTz���ϲ�s���L)��V��b��:�m���2[dX=�%?�I�M���^j(�����kK7�5�9����][�1�G@��M�j��I���d�����.���Z�ۂ��:�U�:+++���$+�����7��B�=D��� j��\_T��qW�c��V��O����p��`1�b �a�I��^0�=��ȢP��[Ղ�&L�I0�5%^ǵ��7�~��%�!1An3R���`��vA	h'4�@�L��A�|PSOrC8�^��h��07���iu��`�`ܑ�LxAgҗѷ��J�`���ҁ��oϚe��"��E��%Z<z;�Su��<�0߷����9
&�m�=�S{Uh04(xW{W�-�k�U���v�CGS���E��~zn=˰w� Q�w}*��Q�������
��eTO"](X��@�`N���?��bN؞Y<��.3���٢w~t�q��7]����)�Y�h��l8_t�A��N�?[L����ڂɦ����K\�a �-���g�@�CR�[/|�1TC�3��bAae����ˊP;::�y �T��,�qu�&Y/���n�uyC�7V'c ���-^X ���ń�`�f��`3���3S�E$�X��j�c�z����e�j�۷"�T)�i���L�aN+�H���$���E��z�4�ʦ��9����mF���G��`!S�f�����Q܎��_���=di�}V"�P|��B����o1���	����`9W>�ss��1�]J
�c��dBL��x�O���t~���Ѝ�3���c�8lQ1cj~�Qzd$nL/�$DBJ����'�@oQgΞ@z����:�&��_hh[@$:�s#�v��?��/���n�-҄a���E�(y`�kQ��L\`T���6�/�:R�ܘr�����F�8n�QH�'bޭwn�A�6���7�����	��y����)�蛚r>��!<Su��uZ��@����B�JCK��ލ�����)���1aD���7�`��"�G f����Y�}�̊i��VV����`?�8^q�hw4 �Gc��}bh+=�����Ӿg��7�@9ޖ���-,("�8��-��
*?7����`s��MF��Aa�u�bkӑ�8�r3�Ss��(~ m{{A@�ʔ0�+�FX��sp��J�s]����q[b6���*�p
ӣ�%oB�N�#�>e�u�����Mq
1hԱH����3vqG�������j>���~GE֦�4���+'�	SfNNzr;������B��ނUP�����
�|!	� %������c�� Z�P�����C+Js�����"���-��in�'�m ��뾈�^�i,�7�&�B�6�މ�|��b����n�l7$f�O�	L�
4lpp0A�����^�8��	y���G�4�LD�3�)��Dm�#������C£84)ݍO�:�����_�gKF�Vzy���Z�ݽ2L���Dg�ـ$$�����S�����L9@}^,�>�}D�A
� {#��P��ܝe�%���z�IP�;%�uza.I#����,FA����[��$koF���1�K5(
4%'�����(�֢pp?�.i�o|�V$�UE�	HjR�_�p2��r`���]@�-�346��)�wuuE���䡥������XѴ_�5�ݼ~G�9x��|�|Ԓ�N��%s��|A(B��ZQP�&�]�+*
p��x��H�x�E#a ��(񥗠�A��̘A�.� ����h_ƴ=�SOwC���#Z�0��B�!��V�-��ZC"*��^�03`^x���޻��{_�sy��sg��6���PЮ�**��=F�����<$1�@x����&g�R�����D��A�:땶�w�G��X���p�&�̰�8R^3҈3�AAڶ���&=��������Tl�md ��9��NdOLL�n��7�Uc/Csä?]�x�B�-�\2?�G/ds�r���Ɣ����]��&$�/ɛ赌���������j�?4�>c�!�R
 ���b����:��ZrӁ��-�~J���U`ܝx�Yh���=_�T&�]�mA�>������$ㄟ*�UȰ���dn�"��Lp@��i��--KC�7o�D/>�&�������;�������S��cbb�^�����(��			K=O�E8�ߞ�V�*#����;�V^��GS:�K�-��-YU�]���]7�N��|{}���QVzU�#�~8~��D�2f���#�q���<Ӯ�/:���VKb�]�wN��J#O^��9�R��(u�)���8�f�j���d��1k�������&IO\��+HxC1X���|�lZ^�×U� O����YJ�V��~%!f����!s����u�?>nxv9R�wJ��<5$4�a�B�HFr�q"�㈗_��'͹�����<�#,l�ů_F��󧂌���J�_^�����mV�^�����)l7��Y��	�:%����2��#��;�Q,-��AC}}�9E���R���s�D���(:�����F����������. �X�y;;�.��E�(��� &�����9����� 8E���0+����[�>���hh4��}Tk���C�!,��9sm���T&1���<��I�}����+`��>'\�!���9���w�X��X$�e�������2oE0 &��e+(;���8G�=��P�F�al�ii�
���Y�ZM˙�9��Q�G�����Ճ�SZ?�C����w+++���#|]YYId����Pv>��R:��\"�� cmGG���̔��_500�Vp!nnn�� ����o�d6�p���b@�<���>��k-	b'"���*Vy�s����&�r�h���ݻZ��-�RS͕�냥ġ�E��K���e=-�$<����J:ndd}��r.!_\�ܐ�f$<��(uV[����<�r���b����~N�mX�	�?������/±��ۥ�����t�w�@U� V>�~R{���{��ͳy��0�R�`Y�7����[>��Z�E����r��
'�ko����,������Þ�4�,**��"L���3_��냙�<�4f��`�e萷8:�þ|�^�L{���p���p{�T�պf?�����c0��g�.������f�ıCE�o�n���T���fA�<�^��$K,�'���|^[�3�� j�`�[gfR��
D�WF����w��
���=�,y�����]���(aSuk��A�0����B��������8���5��H�����}2��q�Q�⁁���X(�R�F3�����H��066V`�J�ipSc�>�H�mu,B�������l�Ν;<�����onEɃ��x����ZJ��T����zz�.(f�j�-_e|���(�$o��ڍ(?Q�jik���K۪[I�����h&$�����`b�0��>�ty�|g��٥���7��N�WC�A���::�~85�iMi1�)�3=���X��r��X�����Ăg�I�=�{�;V<��c"���xx��3Z���Y��\�P}##�}�ϒ�k�8���LcŬPeUKh%Ði{[ٜM���X�n�3G`Q
�����_�lJ'Q�����|��.W����Y��b\F���b,��=eF&&�S��7i����V|,GXQ<�g���jJ'��gS���/�cYH���l��'���se8��
�	M��Lz"�;t*͆h�1M,.�rHH�~l'���{�?��!���ĳdگ�����x���KJ����#ƬY;f9B�4�/�7�hVh�"��?6�R���5�[���v�r�dJPv��]-��{����n�Y���Fo�f�O��E�[����
��χv�L��Q��v���6�y�7�j�R�9gBt���H����y�`��U�Mglk�>��턺Ї�7�� n]r>_��rHܢ�����j�E�;�}p��풀@\U�L���c�(7��;q��-3RlON"t�+�(2Kz+(3��sT?�߳9�B�q?��ˋ8W��i���tK❺�f�S6G��o�'�&Jy|����~RZ��1oIW��t\�}��ʧ���$�^���,$<[�l��*I(���+�1q��GM� �1�������
�Xa��={��+> @��̛��֋�x��xE�������QKX�f�5����8"3]9�)�7�5|�'���K�^����w�ry�����27�K�=ε�Z�h,3�z�K��#��ŧ�Y.5EMA�Cu�v��b�0�ЍL�ɯ]*�r#B�DU���$4��4v�x��rE]HO���Y��Ve��U˝����T�Occ�������P����d�Q�q�A�h醸Q�gƆ���#����2`-�B�����uu/�sV�a\�+�z^=%����~�\PŌ��n��%��O�J(3!������M�~`���m0���*-}v�ϝ�l�q<#�w~nn���xbe�p�imq�O��I3aAA�fK�������QQ%͗232(���C�1�HK{��ff����R��Y!�+�UB�B� �Z:b�j������}}}�P�f1�~3i@����y[;_&%-M�������sO����{���n#���
<?�A�C���&Y��h�14�F��$c�,~~���g�d�x�ӉB���^�G��ѽ���<�~�E'?�dd<����_�6�w�����3B�wI1</��-�o�$}����'�aY�����a� ��.�3"�j������!!\"�V�-3+r����dv� d�N����E:�cUmKƅ h\j����)]���А��DOu���XM>2M{�\qqq)�s���?_#gR0Q-�me�t�y>~������%�j�Qo���7�5M���O��0d��� �ߖW{-��Op�N�0��HMMͱWic?�I7��Lח}�ʘ�(wn,���7l'�	}!Ng:�q5-9�� +o��e��_~����~��Pu}[[��I3�y�t�X�(� ��|E+��e#��-H��2�q��!!3a:��`_�J������ᣚ�������ZFj211Es˝;
E�wY��ExJHT�R�Z�H|�Qgć$]=��k����3t��O��J�s/CU�c�>|+[����d�b���0R))o����y]���̓` 𡤤��I~�y�{QЛ=�b<��l7�`�끽�j��8�sxCo���;���W�����*��c?�0|?lÚ��-�ܪ�lho��;� Kl�c6��V��o��_�43��:��
���ǧ�'��K��	���{/ji��T���MN�n�z\}О�A����v���%z���=���1�%?ٝl$.����%�-�$%�ؒ�\Z�tc��=�ٌWIJK+^ĺ<�iɰ������^ ����=)�C��SU��!�#�~' "�Bt�14wt�U�=��{��=܊����E��b,_mQz���x[=�,*���'�5��5�헬S��gz�k��\��Z�O�o*��L����(�1>Cup�	�Z��su�2��*jj�Y�.��l���c^?��~�.VGS���I�s��]S:$D���1�P��{��q��o�C��c9�E�"TTU�u����$j� Ny��O�R*���c���bUkfr2���LHUQ���Y�-������X�� �ђ�6�h�,ls[9�X
uuu���.�v5]Y-p[�<ǋ#Ɛ����PQV�[��a��ߗ��i��6WW:p� !�&p��򰔙J�D��7�A`s�92�XA���ܯ� Ì�bqw��>����FNN>Z�:��s-�eb�y���WC�z�y�n&�
!ޖ��2��G|�5��F���R�&� ۗ�B��AvQ�6�h5�<z�訷8�a�A��1av���v����(��N���u��0�[�W�[��:��G\������=T��X����3g`b/@w BS�a	�G�={�bgɑ���N\�^4����qk��F9j�2vG��lI/�:�ى���3� Rd��樨�7�;�����-����n �PU����Y�9��D�7�
S���g?��1��wR�  ���|�I�,��]?G�'�{̾�O�����W�%*���s�/~�˦w�м�̃3��Z��kM��~|$l0�k�n͐����	���j�1�.]�,3S	�`=::����Kz;6!A:|��y.�ı��+�a62k��H�],&-�+�����D�6���q���>����w|��ʲM��SO��W%4f;��S&$�d�L8�����d}�`|�yv~�n��E�z���5�|+^ �g}6�:�G�
���=�sUG�4�V����qT�dFr��y`� �qxlZ��y\��RA��u�1S�6G�Ջr�����i�ή�WՂ��9��'��7_L�B֗\	����m\��􌌐�i�仯*�02*�����#W'59
�R Rï��%�pB�/��Ƹ}�0s�on�6\5�>d&R!F&��Hl�]�/鞃Zos�x�u!ܸ�o�?��x�Z��̥���ӳ�C�p�L��m�5�+�SDY�F�%�V�nt�^\�&�7��*�S����It�� ��3l����0�7�yp0u�ǏPF+�uD�R�S���6�ӻ��_�g9�](E"�� N���K�(�QW����J���<oE������
Ik���CGSf
V����P�ƶ���w������q�y�����*~���J��kkyH���\�f�f�<X���p2|ߵr�V��×��4t|����6@O��B.�`�=�'�؆A#��BTM�	vԱ�{h�|�^t���Y!#C�!@HPٷ؛���>��>���Y�Uy`ֶ����R�p�\8W �dӊ�/.�}O����1�w��u��A��ǽ(�Ӻ�~ԡLZ���`w�~�|�7�G�$P��pݙ.\��v�Ú���� z�6@���?;��-��(�� ��*?���Y��l�8]p[H���P^^~�مG�� R�����'����Qt:==J���@�wɨ�؊��賎?hʁ�>�wH��7��ihQ��`��U b���7N��I.��
�
��x���z1����1冚BIӱ�b�L9>>Pﶬ�/		IC}�;�Z�C.��]P;���'�[|����?�Pt���6w�^h�7Y��4��J��@aP?iE�42���f������94�����"C$s̫����5�P�=��õ�T^e�c�6�s�IBd���:멃H�(��ݶ��\m�#,Ec[��f��|;">�f��haUO��<e:ؤ�A��n�٭��D�����jV��<ƹ�p~Tj�oI>���d#�xЇA[`/T� �vTS ͜>\=un��=�{e�L��n�}�ؿ��fd,�?���^�% �t���t����R��>�@��Zu��a�=�>�||��~�~ݹ%�Q=�������kk �ޞq����G��\� ]4Jq���>~�f� m����1�e>q���4.���$�%A�/;���-�(9�+Y"�F���Wv��ǿ����T��T�v���'��!��Q����ʨ=��EU��a:��aYg�)l�� |A��~�晓�c��SUEE*��P�hn�#%m�_��+�H�`"��ӬPĽjW�)��݃q����iA�x�%JF�g�
?16.�z�
�W*��_`AD�97�f�fte�5��nq+��4��>��{־8Ϊ�cs��;x� �(a�*+��LC�����(��L�Mx(CCG�05�Ǯkl�w�p^+s�� b��ydhbb �|iee%j798D4u���<N�\���ڔ�Z�^N	g	"y��2��V�$�8:2���/G�;\?�r������䍐���J]�\��JKPDS�=H���ttb�����+����A���H��V�RQ��V��32x�ϷD)��i�X\��������	���t��:���q����4�,33�7#9��F�j��>B�e�g�&��[lj�3?77��xϾ�扣,�_��4X���

D�+4�j�IH�h�#Ӳk�;Ah�!���e}PD4��
'�����y�"�GD$��K�^�bOG��J�����%���9p|�8Ey�4|]�j�c����b���[3,��K���z�������ߔ��M�{�����3����~�)��gc��隙��C��n����-� ;��:�;_��t�{�'���X����Yɶ��|�Mgg�ys�8EH=kh%N&��>��]��Z�$OG��ȧo߾��6-p�)����哖�� F����~Ձ���F��x����,������}u�6����ҫL�r���@`��0񸆍���K@�����v�2�r
`��ǈKHX�-���uu!������Y��<�@Nb���I�.y�ß4���1I��¡q8�ؔ���@ZP#f�t��d�ț����T*F�W��~ffƈ�ɪ�����R��"�'��E�I0KKY�C`�94��3�OA#
�ң
<T_z����F󬭭G���FFF�4������ai�gb] [?����ly���8���|���D��b�n����\�ڐ,�a�����{6��WU�&>F6�QlƧ�A��Z�S����J�rq�IF`i��h���������}�ͩ �vA��A3 h419`YX���Ң�x�%i�ezJ�Y{ُ�Gv��u�u��q���4�}�MMM��u״C?}'jp�E���68m�LzON�OH���F VUU���N����r�΅WO�d\h����$.���\12<&�L2�|�x��9�ү��ik�
iȻ�R��������~��O�������8��k���ݸ:l�fAf�V��@w<M#�ZF���$$ܰ���MM�Zu��6F��Wd�Ӓ�z��LmN�������l�hs�Y�ǫ�LO����ұ����]��c�+W��ɷ��%�=����E�:,�,V���?1��n�UoH���y�з8����O�������R0k%!!qe�����A�ḻl`@���
b$rҡ�IG��bvu\TT��~�/uuu����ڻ'��h0!�~��aJ/`r�Xz?u�fJi��F�it�̇���`��z��z�����z���Y+�q'�f����$]@�(J��V����@{�������S��[}Ǵ�֦˲9M�ą������h���M�:##C��Q�8D�g�v!c4�b��(��S��������'�Y�W�G�L4kj:禧�)s���p�l?��gI�'c /����Bh��lR�D�� >���*jjBI}>�Ze��,r�[3@f��A^�L	����]hf.q�{����걖#�6L6��LY}�|�PW��.rB�k�-	r�\Xe�~�嘀S�)�0E� k����-ӳ�����1ܸ��22ζg���t0���"V�㰇����'O� �&�Wy���nl8�L�>=p���ňµ�BE4� ~�H�ݭ������Ϛ�v&��m��}���N� �AE����3�>}cy��.��W n���r�/G�p��s������i�N���7^o��E0Q��M--w��+��$��}U1��Ū<�姃��7(�(nj�W�����h_���-	�~�*��lh��,����� Ɂh\��x���3QM�CKg@�31.��lL�v��Ӥk��NG�>1&%����>_i(�R0��D����c�l��E�S�%me&�㝌�{Xb��u
� '���ƙ/�7iL,�&�ھ���˅�m�s��M�)���9Ki�ugc�˛��I��v���O�#<����MXA�B���8�c`v��Z�2Ѓ�͏������ݛ�ݩ��Ȟښ��q�r��呋���]	_���X��?�/k���)3��(��:������K��(�W�]޴Z�=�š����/*��%~���4:ON�}5�:G��{�W=x��-��t���Js��R1E�bb�kIN��Ϊ��p��{��R��+���xn����t7+��)��:�9B��C�iA�ZN��Iթ��̙��#C�R�y�������ЩE`�ȍ�±�b���u��/|��e���o�W�Z�C)�;X0�J_�  5�� �Y`�~�3$4Tz������h��&K �x�of�UV�L;s�% 5r]�}hd��B=�]�n�"b��ě����^�2{\>XO�/�p�/?������U����m���LV�] MEG�7XfZ]$\i{h�'|~qq1��V�H\2k:;��*�R�E*��C����ݬ�L����$	�x���_I��$VT����Sʠ.�}��E׾�6�����=ˤ�b�D�`�=�5|/�+���1�L�I�[y��/��~��(9qqq�>��aVIN����q��gϞͭn��t-�8/9~��)�[X�_{?�;)��`�A���­@&R��7G���]D~�P1��d��c���j��xᝐ�d*4�3DQ�FCJ�y�H�Y�n��K���hB�'�Y�iB��V��Y�J��.=��ο�:�9���^��Z�Y���=��ֳ�=��{�+�ӢEV����v���5h�::o";���^->&�d N���(���i`9L��?$"�W1�궏a����e�p�2����cv���N�����A�d����eG sl۶m<�yB�m$%�RF�1~~���N��iݘ��^�N���6�6�����Qm�~� 3"U+KK}��Cɜ^�|�wl�2-���
��n�_sm5�+R}~?ȭ]a;M���խjo���fXW��D[A!�� L^����✚o��C��1�Twg�h)��F���x�cn�ea3��V�ͫ�@�VS�=W�1[�6�(%Zn"V_V/�K�򼛛>T�ϕO��+v��!������י�������Q]�n�|�6H�Fz������|R2�x���2�v�{&����ì��/[��˫ԥ�ye�W�F����Tl����/_�/fa9�A��ݗu��X�=���@�� /�`|L䤕+Vt�F�}�m2[t����П�����!Oӷ�^��T��[�04���-U d'�t��C]�Yx���tR��f�J�)YPc5��@rr �̲]k��������R�ng��{�3г���H���]g%+���S�{�u�j���˭k��]]���
�9h���Z��~�E����P��~����$~���w^$RW[��������Bo�Ϗ��Mǖ�^2[��D�����?��u(�ſ��233���}��-fƓg��O�ך��>�����k�j�|�{��}zTz� �s5�U��?,����W��N���ލo���{{V-	R�q,Z1��P�DD1��B�T�#��܍Lc��:���+<�r~Oˏ������'O8�
p�y�n�֛fK����Ր>ׂ饾}T~�< h�@���C�� }3O�)z&�q��А���t�2H��7c�x���~��x%~�b����YR2��G�o՗I�F�˺�B��S^��`W��y��y���䏐�t�SP55�L�v�.�1~�-2 ����5�e9�YR��J�*�|G��l�6�Ns@MX����Ǫ�Ĭ�J����t������t�LR}�uѳ[�����,���l�	��@1ǽ����J�>FEw%V>���GZz:��C�E��8 ~�-�4褗����ֶR�_��nT��h���UE w���]��C?�!v>�n�d�C�k����z��s[��1Qo�<�5��_�	(*.����1V�t���k��FD�����O%j�/�@�K4f|||T
A���6��/�Q�XQud�\������
���n����@��-�IH$�%8�!*�9�uq�?A�u��	4��ޅ�S�$C�.�_YI]��g��gQ�@�r��
�PV��{M5�Q0�1��!I7�NI�RɃ�6�<�x��Zvvv�/���}�C�����QTTԣӑ������^/�7V���T��*J�ض�O|f#b�Zy�X���Ǡ��l�-�uu�ϕ� U��1����lr|�%ϽG��*9�����p/��}x�T�����>���Xy�&�h���l]Pv�\��#/^SZ�@Y�~�+d���t��0ק�Ŭ�[�8B��f͚5�����1�9�w~������Į��a`�i�*�3>%*3��~��Ԃ��4��*�"�MM�C��#TK�S�k�轭n�����\��U��J�.�jP,�����h�։V�ǿW�k����sr������f�̋-^[�>8%���f���D�V���!��_�O+**Z�b1����>�Q��_����g���v�C�~CƊN�_!Xn�����Y��uTħ�R��6�{��,�11뇃< Ӈ�QBq�q�{������X�<=#A��錭��!��#6�t����]>Y�4���W8Q�^	Y�E7���}���h��4L�P5�O�$�Ƞ:�9G��h唋�%nnn0�D"q�3�a��q�l��~�ePYW�L�ʚZ��ѥ?'��Ǎ�	(��z�<���q��b��:!��W���s�b��~�&7-��OnߌMi,פ����p��aze�U�.��¡L�	M#��F����c\��3��4X̽�Ƶ�.����V��K_��ж��w��&��{Oʏ�ܸq�WH�`ҟBϏ��|�����/���R�Fs�)�����r�	k��N�x�.�ĖKL "�F..��6q:,��z8��v:�Q��j$u��W^VG���t�D�}}^���܉k "��j7�?���ac�n~kz$�Y a\��Ũ�N��M8���%}�"�<�Sh��{�)m=@�κ��)��ҥ�k<�C�^�*fG���jV�����-�9@�E����Hス���ǏAm����Pz���Jn���#A�۸iSJ��j�i�Mר�h�d��|���e333Ә)����l�t1wN�w"�a�b~�g�t��|����ml,���~�4�KxB�m�-�ߵ��$~���c?��������=��|T����J���b�}�>�C�9� YR�k�*H��
���g'#����աq�.$���W�x,�VRR2�i���]5���u�t"�ENm�V��4�����g��p�Ѧ�"���8�)Z�B��ӛ�>��?�.��f��:���:�O���)�Sh/���=�����|����1�
�A(Gs�����zgQ���^ul�,9�n�~�0�������B��Ç����l���4����*n1{��C w���g�
÷��]�v�*���*�~|�

"�km�N�u��=Ŝ��,t$*�������,s��kEa	��O�v�:+�$m��o�}���ѱ�{����;��]�Gw<W���C��mrIގ66��Y��=i��:�H0�P<:s��`��dS&��N��ڨ�?1q���;��4�B=[���˗c�8�0I�"���nڅdY��q����Έ'O6@�������]vko�e�R@�I���*(�7�Q\^o}&���.�����H�S�5��Y(�])�}5L�iP���]��#;�w�ccբ7�~�Dgg��M�D_�h����RHTsg@�|Z�WE	 �!�"P"��\�vM0*H����6�F�_�<�o$���E�P�qM,���
*��+����&)�+�W�Y��U�F.�l��P|���T�[�FG�!oٰ���*���XdMŁce�WXL�
��``FT�f����Z�%��X\Q�_�8�Y@�Dhҿ�;i�5�	����Í�w��RE}�$K�0���Ϸ��ٛ�::��>�YI%B|�=��ܶ��0��&�7S�C��Ϫ��D~Z��8�,~�,����ɡ��R�hNʽ�:Ff�s
E#1)��]NZ�fJ���f0-������Z�xr�ӧ
L^�C��qt\�s.$w���� s����,�p�m�{g>Pu��صV��eܒ����4%�q<�t���^��EU�gve�������l��-����q�YN||�5#��O�[[/�5��
����m�\3n��_Մ:
27�|�����H�6.V� ���Q��e��F�u���0`�6&����಍1I������j$R�=nq���nxt��Kv*�kjjR/t�6bvoF/}��B�x9""���/j���|���R�:@G|L�]T���V 4X���<�t��#E�OZ��}� [__��[�wS 1������Ȏ
H8�3�65���:uwPYt�����t�BtC��kb��3{$���b��W�f�s\�,���&'#�M?����h=��[r_gō��2=lܾ����ﴒΓyw�.7��x߳zs����<��O����ٹ��'�f���_k�2�z�ȓ���q_>�:}�כKm��ٍ�ο/�l+5K��� &M�A/�v�e��Z�}�B�!�~o��5�ͬ�=;���E�t	ޮ��6T�O6Bexb��8���WUt�W]�b�ϟ?��탿C3�&�!.�{r/�K7H�H6̻g�H��XTL��\�0�1�hYhX�lt՝���b0/��ab����mTӼNO$�6��;�o<lڴI�wɛ���֢>?��R�&�������g�����5݃#���~ű�zw��*憫Q�<�����U  ���M����7�GR��7䲠��5��+ ٸ���o�+V���%C~<���DhI۸b�`��4��ArG,���f?����e��A'.�uX�;�=S=�������~d�P81��60 �$��<^�a5W�<V�5wV�%���g�n����b�Թ�"��^���G%�:��vH�A��W�o�� �.4���͛��Մ"��+۶�7�jI�����s�>� ���녚�����$W�U0=��F������{��N7\�1KEo����Rv0�� 0�\��Ӫ*M%�Ƣ\Qā��y�~��'�7����B,����v.Xk����j���F+�$��4y���BM��C������hD}oT����Xxcd؜2������孅�����������d��u�'�0������w�SbEm6�#5Q�r��g$�\�$ �_��X(27��'�Ӷ�l��1)f�ak"�{� �[9Ւ(0	��&��-4���M�����8��$\�i!/�9��:8:��? -zخ����yy�����������{5�_�*Iz�4<5ԭi'�fҤ�zC� ̈́B� �s5�e��C�o�C&����?�oMp�/J��-�2�Yfә��y���u+�����ՎX4�E���k����u����q5�AېQ�ɬ���<��e�MB�x��5ˍ�L����QuJ+�����%�o�OV�r7�n�4_@hX{"+;��g.^^���{�J�宵����6��U�����o�h�;�p�%i�� |`��r���Lw�<!.Vko�ת|�l��7%���N\\�4S2����@ݠ�X�|��6 �<f�k��3�%=%l�NzOH�e̴���HMZ�M�7�d���o�k�:�y�ff��=�e[��M�M:%iL���'m����$3C!��j���ߔ�G��4/����LP*&��#[�L[�|�� �u�U�;��{	B�0U?�iQ!��o�%�v�!�I#���C��=��O1������z999d ��V#�:�>I4�s^�о#a��Gž�<�Q�jo�#�B�D���ߎC\�m�x-tE�����"�����F��l��5ݑa��9�sG�V!e���헃�
[!����'HȅN���H����&���ڮ�v���P��TI=W��ۜ����$0���2���O��O��	���Aw��Z��m��Wq��s�F����*�!
���OW)	9gut�NR)�N4�ƊŞ�DpHXX�]��B��,�Ѵ��g̢�R'�$z�]d�z��qZ7��ll��1�������6��_� �p;v������t�fټf���>� I�9� ��Zvc��NـK��m�cŤ���=B�V,��-�'����߿���F߿Q��p3z�����|�351�hDI���ېEYXXl�]�J>�
>H௩L޽Y,e�����o�����ϛ�jo� �>�^��F�m���ݖ���h1X�䇢��4���2.��yr�ѴHک�|!�V�K�EFFV��<�tjj����WΏ��UyB�m�v//��h�������{'�"?��^�fS&靘��h�u���8�X�����ޓ����P��b�E�	;�~��� ����t��
to}	B���ӏW������_e>��G���A|m?�;��al�R��OK^��#1�~A��e����4_�$�='AX`�K3�$x�b�\��#q��3��=t ��
�������$�
�&ל��;t6�x��$t�%��ˣ{�Sp�h���>���% �?(s-�ԽbJ�L��q6\
�[/���*���H���*�hs<w�T�2�ߦ���e�"�����h�֢
��Z߹������/�t#;�˙��9��!���4�c=���if��}���c=}}E!�Z� ZH��mn��!Q��[��OQU�3w>$.���2s��XrTV� ���zo$��p%Y w�@��� �:�����f��=1118�g���i�/�il�T����D�n-m �>�N9��X�B2��ja[��"L�����%�J���O��\�����D䱁'`��Ā���/�{�b��v(?A�N#=:��h�ק-����қ���~��A���r�g��2%o��ܹ}e���tw	@��$H��s):���X��N��HKKS�Xв"�Z���*��I΁YP){����c7�y�c��D�����pby�ZrM!��=��� ߈Y���+�����F��Yc������2����@��������6/^���[����0�����9]\\^ggo�k�4�	&PUU��B��\7>���H�e�O!?<`�z��P��@h8=�.�lQ_�eCI:   �>��3�?p�^��v���雒r�7�O����`}���#@��\~~�S;#��橲���=(�!��8��
�%�w���{���S���$�w���;��;� @��O �u���ޮ��E���%� ������w]�zn���$'��#�h�]�Ҕڜ~�w�~�.@R<9���#P�Ԡj 4�yidd�U����Ք��j`��>A��[��AF�#j�!��C8L���*p%栍�a����w]�	� $F7�E����<�����Z(�`�U�fA��I�cp	���g;`�ɗ9r�|D�_/]�͜���H��RQGJDM:p/7�E�L���ӎ�v���Q�Ǖ(#��_�^F��|4V���C��y~�GHL���������;��]�=:���� �ֲ`�J�t�و�q��iH�M͏0f��"�7��E@�i�����aB(ף[��F�ggg�NIiSw�H~D�@��#w���'~3KE�p���X��#*@TK!%�5���!�T^F_f@��@&������,�ѯś�?�#D
�Ի
�84n6�#�IW���yHYzTy�+��
�Κ 2ˀg�JJ����D��u���@���r��\cJ��=߅�|SLR6�K�::���k�M�2�3��m��Ex��,u>H��@����@ ����T+��E�(f��t�������@�0׀oxX]�[-�V}���
K�6 ��+Qso�����E�Y���������fS�����U
i D�p��I~l.P�>�:V��\����t�[G�#��lZ�.̈́8�>����F�H7�8�$%M� ^������q�v�q��֓t�*I��*�<#@֐������n�K���Hˍ^�O�k ��W�R�fl�X&:��'������ad�]Uѯ32��_P�L6�ŷ�VVň����V�֜P,�eKǥQ��P�
ڛ��kH�sD I)\ʗ�L� ���n���S��߹[��n ��y|p22Ǘ�ߺit�u�7%K&:��\E�[vVn��R� ^ �|��ƿ���C��==�WzE�W!넄�>��1�V:���p��U:e
��O�i$ҿ���Ħ�êw��}�l-T���1�5f�K
�N1��zR�u��$==-]��d@=2�XI�!<<�f�./C��!���q�\�&�i�l6�������5��7�t��������_U�������\� $�E�<�]���"�<������t�廬d!�B��Uϡ��=(_Ƀ��^�'B�)��ucTkƯ�zݿ�.Giv0�Y	�--��`��F<�u`@Ŏ��p�F��^��BAY/L�y5J�|��-�x@���۵(�itH�c��Y+DPd�`F��Q�����q$�ҽ�%�c�h�&77���l$�)3�@��<���mX�=�	��sXpɐ�(��q�&����ۣbmpl��Dt�LdY�4Ru������:��)H���B���$���S 3��_(��Ӄ@/���$�ƅ�}�������MdQ2uuu�zrss��W>UA��V��'��s��ZL��_�ta�#�𽍖"����� ӏ���;{���Т_Z�z����L�i��������z�p�D{�ʻ�A��*Fx�/i[:i@��PՋX@�ԺLaj�f�A���ڌM��5� y����kz��~1vv�҈�f�R9����Li���+}j{�zbں5d�U��U~� P*d��VB���<$S��sj�|���r?@3���^����Ѹ��*:�����oL�h4��Ż�v����s\[O�U�"�u/��mP����/?�[(�$Z�����mT}�&�`%�T��e%��k0��Ç/XX����./�<$��$�M�':�P�zMl.m�M�F�В]˦PP*�
!�|/6cK����9Y��Z���'�6�'
�H�Kx6�~�ƿ>B5V�
�,�S��N\��zz��b��S�NA��������m��R,dK��h݉�D����3�\'�*�̱�q�y�[�Ys1�Q�A�(��8�C�jM۶��`oOK�t�re���c�]=��/�ӈ��6����c���9[jB����������Q��Zooo��,� ���'���(�Y�N�\1�Q�>�}�a�aE����C�Pa`1����X�r@5����Pg����m�C�9|Q4
���NCCw��!p��O�|뺶��MuU����V��]s�E�B�օPf�����WiƝ*�p�9�P�c����Pۻw/���Θ�������:G'*�iR��' �_�H ��L=�y��ә~
���z�ȏG�c�˰���2Ʉ�X�����󮀇 Ę��y��5��=$$� �����d-5QT�t;d���64����/��W@EĬ�e�M�6�'��9D�� �4Z�ԛ>�Ґ��ⶒW� �9��}����T@O�}R�����҅[����PG�S�w5��:��
��@��yANW�(��sp2����_��Z�	���4��
Ҏ�԰���;��37o��տ|�r�$��iG�n>0�}/@��$q�3	����Y�b~��Ŵ@��.���s���(��z��2��(��םṞ즡O�t/;�z���ʌ��}��95ONN����%�g�i��xH���$��t�4�����F_w����+��ď�y���OG&u����{�v��#[lA�`��QH�NÝ*��a�vV%Kq�Y��i�S��Y0�����pat *�rDq�66*l!�?�so�
�E&*x��;��èbho33=�?M��VA��ϠSȼy�" N��::��$5�Ԏ�L��hAC!aax��������
-�))�z��������VQ' 2���3�)�.���n��}Tcע/�@U���)��"�>h��0��w�m��l��}l��'�X��U����DQ@׀�燺��~f�� ͷA|E��u^�Իz�\�A9�@{ie!���^�9g!�F��-���N��V���m�����Pe�/נ?�EݧŪ $�
�h��o��Ѧ	�}[[�6-GA1e�Ж�7`����%�y�oDA4�J�܏J~��֡r�w��`�eAw�n�U��c�aO7��<H3Rh+
���$:�y�R? &HۈŹ�[���%��o��������C��h�җ��1��#	&z��h=L$-=�D���h&���Uu���9�!��բ
| |BϢ����������	�DM$C��qdn �3�M������+ShfP9i(J�l)������:����V�� ����𑲵��E2��xI���"�%�=��=��
��h��F��NII� ?��R~d�ٷ��[�r�Κ-��o[A���wݻ6l|���F�'1 �C5Z�S�6���NJ(Ix���px��+�6 %��_�~@�D��\"*���p�P�#�DA�~��̙3q����� �$�����Bݺ��V���`K ��� v� 7!�@?��}��IE���9#}�w��&d��Dx���@�/�w�}Z}�s�4l��!g�d���
=�C����γ�o�:m=�w>��}���`] \Q�z�"�� �@��
)�x�PA��-.ix�[�e�7�vȂ��s�� �����f���W���D����^DU[2-Oח��P�N�u���ٰ53�Dr���9h��6�_oq�ҽ
�/��;��Яs!G0x���iՒ�o������8��Z`��|XG`�[��+���Y�*v�*Fw�
,���m+����vvB����y�o~��l���$Rds!���
zO[-��W���&%GC" �!W���0Lu�F@��UY@��G��s����RT݃� �A� `A+ kNHN����`5��C`F[:���蘪	���`zE}�2y�������ޤ�K��������ab�A�Z�]ꍾ:ea��;-+k�4
|�m]�ȥ/R\�jq�2d����U�o�
�,T�� �DD�w��Ǡ0)�l�i�s��R	aL��i �/GNf��Y���hi���M~ŕ�U]�#��s�=����^[����P})PG|||���е�%���4A���谿���A/L��ҧ{n��� [��V���V2�oiu`c�@�[�%L�DFtA��\ 3h��H����}�>���~������6�mk�~�<�=�P��}���y���>�6���V�E��[�[9^ۥ|�l��X�~��haa!:������`���v5�b���`�ԃ� �4_-4�2���YX��W�Ջ����b@�M��!��T0`h*�c����㗟�[O��� ��7\���y;1O���X��TU}CCïz��e7?"ɒ�6(	`A��]�/}�xA���p����t5�p�r�>{l2�EŅ���̒t��/��M�h5��m���[����
w��/<��%,��7ȩ��&���=�F�y��������!ˬ½rBd_؇{Va�u܅&�5���fw��3kW"+�|L�:Eu$�Θ�>�3?�Q�Og))Qѱ�~��������͔���O�d����*������M{W�reZX �Μ�9τ����#�y3��M�,�#ˬɜlҦա%����S�h5,�:K���%�����深s�2�3|�h�V����c�(X}����%[Q zG4|M:sz(�;#7���A�8�h�8�]��K���,)�%CP;�1_��F\�8�^�uN�i`U�����!�Jg�:�Ƒ,C$��c$��^Dr5F�
H�. �Ia ��Eǥu0L\g�5��L��%xg���Z�L�4\����wFNM7�z6����K �
��;ܕ w
8��Owb�]
������0�>l���3�[��F���̓r=p�r��I�Ϛe��^��;�L���⦻���`��܋{R=	5p�r?� �I`�6��|�@=xX�ql�z�l��5�����Hr�Sn��-f��'�?�`�Ӡ�r�jue��?���A�Mw����,YƦ������VC�m0�P��П��p���:xă��<�'��I-�V�E��`����$�Q5B̳��k�����5)\P@�z�Y(���@�M'(�{�a̐��&�P#;��@O5��5�.V�F��Ƚ;-Y2��!l�<o�� ���&``���P��}Lj�,6�G7��;��)�}����ܛ�]?�3� ~�0�S��A��NO2�f� ^�d	�Q��1��la܂��:5�Ђ�p�B�Q����Hg;X�#(�I�,�U^"�ryբE_ާ�~yY~������	a�ˍ�'D��ě���n�7���^��bG�����%�7�~1�f�}�x����{��4/�bhc�'�lw�x�����<6݉��>�0�U��Ln#�}м [�aඃ�+>b�k6�d�~�m��}��,X����]�E���Q�o�Q���|�:v�(�K=�gZS��x��Jg.���0�\.���a��;��<Rs�9�`s�	�+�0F�B�� ږ>��C�%����дݡ����]�G��ׁ���8���@��9�3q���v)�tȶ���������J		=0OP�X+ a��9}�h����A�L��=A���ى�<�Q챫e�d�Ŏ8�_Q�I�Q.VL���jN_�7�=��+0�1�1��0#r �y`%6;s���6�[���+�n(ja%�b���0� ��-Xo?PhK��3��XC��8���P."�c*��jw �|�qr0=g��<��D���9Z^�q�8�1�uI�  ɂ� M{� .��b\�(�ԖJl6���<L{=�E�� �3B̯8����A[ڠ���V�A�F�Pg���A�0�!Ѝ��y��`�o�F����EY@:�X<�A*���C��zй�GN�1ȡ��=��������64��M�]n�`����uє7�O���d0�1x<z�P�I!xyV��z��<+-���j��G���!~@n+�ۍ�J��7���6z� <&�=�=���[�<�#��t.m*hT\[�=�6Nw���2kAL(�H�2��[��f�"��K�{Xg��,��)�A+`�3�rK.�� 3L���<��1���$�G�5�&*����a�%
3ʑ0иBἇ�\�t�� ���'���=��@�w�F1�-��߽��y9D���}�fl�ϐ���V��F&�̂�l�R.�}������Л#O�4�ڽ��]柈��-ւ��h�y��	���롣7p��!x,�ėNK;���z���Ή�)����߀��7���o����d�|��,������o�����?Tyß�m�$��q�M7�����W�v�(���(��%�mp���Zv%����.����)��<����1�R�25.����w���x�,�[������w$�R��@X%�����~�O^��v�����*���_ծ�1���#��9���F���,�o��l,Y�x���nof�Ϳ��:���������՛y����d!p�la��"�LK�:�I��v�\SS3���o:{��#:�rqq�`�s��U��\����w�ȴ�`k��+&ѻd��;��`N���І���C��&�ᶌE�mĕ�\W^�m̑'z�Z,�;z����&����f�u�3�8^��4�V�naU7����Q�*e@�1�
/PAGq)�-�w;,Y΁D�p��Jg�]���HB�}��gqcK�NgN��2|;<��eǵi��8g���4���ma�mÿ�o����2$.'����G�a
�Іی?z�ؠ���NÌq��|u��_7 ����m�9���^���#�����q���pM�ΞH����t��vVc�@�hÝ"��m��w:��NK�Nk����V#MK�[�vǷ�:��9������fh�yP~��ݲ�8ۑ%|]�Sja�q��Ƴ������#}a�7�3��mE�V�ZZ$U⒣��n罠��Pb���P �X/���FÃ!G�}�AA�����xP�]�{0�A��G�8	�S�Ծݚ%w< ����H<��=��u�ʊ����ߒ%ȟ�ݲ7�r9��P9T��n��Oa�5�!�ȴ�
.��~\Hp+L�6�nq�G��6�U�� �5@�G#XA&��0"����x���&���cp,���~���ha��Ex� �p���J�����v`j>�
��aj��=(^D�8FG5A��q<m7�m� ���Q$��ë��r���fl�0ƅ ����	�@n�	�����6�{���XW��~8�͒e	Lc�6�9���K���/��w��1�P"���k`���Jc�KnN��cx:� � ��Q__o����]ϴ`��v���?Y�$���q`�3fc-���i`w <�a
{ (�<�Jm���A��_ ,���n�%�e�EϘ��Ā�� �g츶�І�ۂk�!.߇��6D����6"zH�*�6D�w��:=����:��6f�m��D�������w������^_?�Ӕ��ǂ�ҟ0+7箯��y��E��������(�F�1�^� 2; 2��d���5�hǨ��D,�n��q�ȭ���]n����[,YZ$G4a�J"��Vk�� 1�� (�bFM�F�:�?`Ѓ��..lv���`dn�Hel����Գs0�	J=y�/=��a=n�`(�l#N���"�K�vূ�ԭ��у�@����"賥����v=�6(�C����{9@�W��a<A�@�ژ>3�e��(k�G��|sB�������2�B��`S� (9C1�W��NDp5Fp��>�wb���gG]]]C`>�!�%���b�3�][oς�bzр��J�`��w�L����T�
q��U^�D���Qah+��]�U��GU��]L2@O���6;�:���M~�; ��,Y�f����<"��Wɵ�}455���ߴn�q�EG��)�X6fa������bbډ(?��e��چ��xR���� z)y�$P`���*������	j�A��Sy9 ��0����R�|����� �P����c��)*6"h`��I��bn5����*�
� #ڸŚ�q��gv���-���P�ȳX�j|�k[�� s=;���$�`y&�z:,f+���0��5g��C뮑n�����c����%����|J��Rn�W��S�qmm�Xk]��̞fB�ۉ�����؟����F���c8}���|�Q��׌'�e�u���E�r���i�K<�$�Ý"�l���g:��%䌗|��Sd���c���D7C"����_$t�2��z�J�?}dE>�������Є�O2�����2���_���+�ꔈu���?+<
V���4�㿎��u��(ϑ�2��&�F��n5ޚ(�}}�ʢ��ݷ���V���\�S�^�����	��U]e՛(&f�O�}~v�Nv�Ԕ�?v�:^`m��v;d�jSM��#K���G'&���KM�.}�Y�<6�wf=�;@��j3o��?�N2��W�B��蠣�YV����c���7�A������p72�ѡΧU�5P5�ᨤ�&Y�ώ�d�mQg'5��Cՠ�i$��rO��믧����u�	h�E�'��1t�4�fK�R�k�{�>��A{���n�߄PR��$���I�T�W_=/�g�q`�{w�E>�LmB�"Rܙ�?��dN��q�ĭ#S[&������yǑ���\{��ә�C1��_�Y��/̮��aN=���d���=,&�!�a��"$�
�VX�ߜ"ߟҠ�����0q��lE�������h���T
��B�"�������B��_83h�DPVN�?�<�I�[��ş���*9C��Tiq�*T�|�����R�
U�lg`x�ƈX���t�r����x���wP�T�7v��A�aC�c#"����j�_�:TX&��hμs�g�Sf��w@�X#Z�/��ԟ��Z�P�i�y*E�"��k���4L5B���Kz�%�uӷw�7��v�t�,s9��WLE�7)ͺyvq����J�.?=���oi�xs���_?prk��k|��G}��a�
/+�C�ŚV��IDC��wޢk�2��ag�{��?Q1ȑ�����ԩ���mV�Hځ����>:S���'JL���3p�}P�O�?��zvh��l��=��V�Q-([G�a�\�^-ꬦ���u\i�@���-q*�z�2�T�Z����n@S�M�ۂg3��-)uFa�I؍Q��#���@3�pJ՞ZjW�����d�ԭ,���(��4�"�.�(ƻG�Ѷ%��c���,�!�!�9u&k�d�S�'�*�2�R��s/���zn"����Zo�|�d�5;4f���"���db�fMigف��$ܧ���k�f��>�x�?-)����I�y)b�N^���ՠb�㿨��ء��rxF��}*P\�雓�*�^v
��k9CU�.ػ�.�k���1pC�\x��v�eӡ�R��88#$)G(,q�Z$�����z�V�7L(��.���6���&n4�n]3���'�숓9�5rr�oRs(v������X��@���8ůT�%��o&>�S�0��R;�z�!�1�t���ܤ�
U\�a�m'��IԎ8Ǘ�����bQ��L&:��L�RT��_��F^�"n��ݺ��{a����xn�Ȝ�_���V%�N���U(�Dq�հJ������B�k��$��fe$��3x�����cмǌD��m4��Rg��UrS洄s��W�x���]V�$�H��տ�,Խ��&;�j�L¤���J������I�(���g�m�#F�|*�)�)��"��t���T��x�֦u�J�12��<�A�]��<�ϣ`�ie�'��W!�Lt~X���r���[TZ�ckB�ǉ��q�8#��Ó��s��?Qct䘼���JgS4F�8��w��eD��ΉC?�[iB�[tU�M�&>��^�넦Nn�w�7ڀ�o.�k��{{L��I���Pqd*ى�E�HjV��	�7����K,���E�k	�yo�L�mr/�-���Z_�jo�1Ev4�}�3fI���o����s�د��l�zpb7HW��E���eP�+r��z�)Vገ,�/6W�-)�������ɚ��Yo�?��4����(d@o��|�J@,{uo�h)�9�2@Q����ws�M�L�f�(�i3Pg�ӵ?ko��8�5bQȋ���Ϧҕ�Yv�r��HRS���ki�(���g�a  }��Ώ'Y�ޟ�|�ڞ?Ш{��M��X�$����K�����JN,O0P�yK<fok���lG�w���IW7��LH2[�Br�>���0Է?���SY�9�Q�r�VO�,����Z����씬����Ĕ���觢��r�r<�<.>:��T?��\Ú��H�g��2�zL\�yp}_1s�����Dt�K��3 	!5Z<��x���ZO���&��;���ニ:�}+u����1�T�<���/)+f�!"ݯrЎ�>�^��!2+͓�w&N:~DQ��T��)C��k��ҝr��UU�	��`B�wF�C�7yh�H�;�F�+�)�(�q�u�^�Xj��=�휾�L�0�����=����j���I>�xd4�,�)�lL|1����e�^��ߓ(u�����t��?��o�u���4��` ��3�&��b':x���'n
)^J쬾�('+#�]#�iYߦ�\��2:�� B�iTc���Zs��
/E���lg10��})u�a`D�Z�L!�E�J�O�� ���P����J��r�0���%ny�a8]�r���������0L�.+}\��?�c`�a%f��C�F.u�^� G����1Rg��r0v5ҍ	8�D|J��.�� �e`@:S��O�_�`@���������J�q��h�d�.�t�F߁=��=#:���Ga�?Ƶ�s���e��M�bYL����0!�<�R����d ��5�����\�\]�0��)�i��:ԟ�V�Iz���x�*��j���l��	�b`#=:V����g=��j�b��Q���<�~|��{��7�mUթv~ף�2�Ա�r������dz����NM�d@u�����b�Pg���ݓ\nka̾R8ձ(C��<���{��fٷK��� %����bf����K]�t�����qR�S�t2�g ��n�?��w�T�&yA��'m���F�~.��?�Ni�I���K��u�{oˀ��5iyq3:S?fy*f Q�3��U�u��������P�;��ș��Q�nC�72�zs������ݮ�e7��? ��>`W�-i\��:����6���!�7�m�����M��%���5�����c���Z�z��Aׯ��0&W��{���mP�7��]Kŗ�r2 ��rq�q���ͺn6O�̿i���#���l"#�?�g]x�e?���j!���z�VMjV���}#ī�|�^���K*��dEi���_�>8��4��:��`|w���	�K;V怳����(�W1��Qj���´��L�x���G��1"U�7��:�WԽ���ok��NPn&Z&5k4�;&��F�,܆����ɖ�3����rnvS5"Z�A�{�S^�m8�"Gef���.֐NsW2�f���?O\��;�_�`����
��4���F�)�,j�T��ԯ�}�3��a���Ru]���:N}�,�J�0\R�O��8w����1VZZZ.lN5gS��9���Z�=5<�;����;�đ�߇����E����Fø�/������d������s�����[�7���
�%zm��9�F�nJJ���I��T�ʹ�H��{`v��ѽ�\�NB�%�)�rr>2\}(�ִj�&��r5z�յ*��n��E`�O�Z��5N����@���~��ި���D)�)��oY7�j��rF������]��l�xy~�&Y�u�۝�3[�.A�ya��z��B����;[��X5�,�LS5����%5v�j�j�7�[�S�Sv�~ qb���늶�0�=������-w?�}N�p�	��M���2#�w�{��Ӝ݇�� �vt��Q��u��6jd���.��5i��R�6=�
���WIA��K9�YVBd�[�G)�#�(�{9W�UdI��fxh����'�U@b'C(u�R�r��S��,»7x��ʐ'~9:�fg��;����y$����:�oW(�(���yv9���Җ�Gmn/����6jZfZ�����	`�^r�F���̰#�U��v>v����L��Tg��a�MJ��+����I�f!⪄������i�I��bW�7k�c`I�E�C+�<�8�N���c�0^�p$��Ҭ:Ĭa:K��+�O�*3��u�Tza�d�3���)���AS�ī���?�t;Įo��e ;����k���mrl7����AkS���9�_��=71�$�Zu��ඳxBgH�a�)�u��R5�v���U=��[�f�FzY�s39��D|�:�\������X�º�:����q3J��x
�c0WY[{{Zyf���@�.^�¾Q/�O~�JcnW�Y��V�}O火K-�g)���,פ|Y�m�h�s�.�I?��Ԟa����"�2���s��F��w/.)�I��[��C�����B����Yi�m�@0W4�جW�A&�jC���Z�4�v��Û�1�<�D�ב_܆�Lx��*���5q���q���W#8���>_��ܾ�f,�]��G�c<Xte�i���:���5��%o2�X3�%��i*N\�-�%	Qk��;��z%o⽞ +QwD��OΏ'���#��Cuݜ�,�ň��*�JM��iۤ2;nQ��ab'�����x��db��#�������0/I�y��j�X%��q ��˰����K=8����`ͱ�׶�Ę��O����)��P��R��{�N�4�� ۵�ô���i��
�FŞ���"+�<��ˠ�o�o�T;s�N��63L�����J�먓����������"ý ��#o��j2���|L�C��`oo_�' zb�|·���
eѠ(f��n*ԡL�g��e�~2�U|b粰ӗ�9�2���/۫���8'yʱ1��\�꥕��v-ɻC���3_�EY)f�e����=����=����/h���+�Z��b��V�S7���K�gE@�!�"R@A�a	�X�֕Z[AP�%3!��HXԊ�7������|g��=��˽7s��O:j@!WN ��rDb�c�����Ȧ�0G��FI�ٮ��뮁\XBWxu.�L��,ۄm�߅�X�y3��W����_i�׻��ٸ��Y��v+�i;k��gd$O}T%�Ti;�7���]0Wft�O��w�J�5�����ѿUv���S&�nI"ҽӼx;�\����?ȱ�5k�d���C69��cUz���)l��&�f˜���ܥ^غ�*�N[����F�3��v�O�a�V9n�y��y����)����'�ކ�o���](C���m��{Yk{�禗w=ݕ8��n.����-{y����լ�Q��Ӕ����9G�\ࡴR)��G:�t|����e�&D�|�ѝ�;�Q�����.��
�5�YmVP��#�aa��d�֩Y��OSo�5d;�;V)5�cteI�n%���K���낌��C6��{AD;��$#c�_�ƒ~54��m��D���F��Z{��`�*��ȥjiGlXM�*�U����b{�"��	��fs��%������������k�g�+f���K���/���^�j�ϩE����K��s!>�/�/�j݉���k��8^��z�,���]WIxs�:B�q���dt�ő��Oޥ����'�����uȚ7��"��7|�KA�B2Ȗ78Gܲq{�$1C�Į~��8���v�B�u$=�I�<Ų�Q�w�,���gB�6��d�w#��_���re��<H����Ir(Rv+�Nw]}�x
9K�8�N��kJ��e�X}�F�r���*��D�֥x�؇Dڞ*A��s[[��9b�ӹax�б]�B�6-�ZR(3�a%��Ʃ���*{���j���6<��sE�A#���Un7_�k�6�U،����M��y?���|7�WP/�%��j��YD�9�=e�*�ڛ��;�mT�R��&y��F!��\���=O�(��>��q� G1A����Lk�������ӻ�kB���GtVd�_ݖj�B<��IcӇ�<yED�|º���TU���: {0�+�Я*OJ=x�DS��q����,x�m1:���K�<��@�3�x��6m�
9�.M�:7%y��[��-|�z��F���wW�e���%��C�k�ۻ�a���Gy��5�?8�hp)�3W��	��˜�k$��y{�|l9?��=�5�E�!��-ݎ��̎j}��@?���6ͪ]�����y�b2��!x��+/�$E�O�2�z2|Gz���r����{`���<��_1z�nq�/�ڎ�zU��}��������$[�/���������ks��Y�l���L������Ym���ԛĎ��o/�\hd�in��l9������G!b�#����&oN+(�إ#� ���\G���S������)���&�X��6S�LO!�X]�\I�����Ǥ�fo����eP���Й׏��рt>K����r6��t�ذYr?v���NӘ�@�<!�
5�'��+���p�N��^/��C���䌽<��R4� ���/ׁ��Q_�fɪ;y�分V��'�0,�����cǸi�Z�e�q�R]-2m�:�V �7O^ƍ�������<�\��=�K'��6[�_����������L�`t����f0�C��R�j�d��&E��c�o�D./��"=�hl�J��}U��(}��q�X8�xOc���!ٞ�>!M�J�h�N�(0G(�,$�񡬐�J�Z׍C�z|�Lѓ1�� �AY(�I�H�u�,q֥���B�X���m�bR/6�a��hm�k?��C��k�e��������^�7<t[?��uHorU��G�2�(s3D �3�rnpb�q:8ٖ��~wl}����5�c�
�����@�"KQ��P%�/O~��$Q/�w��<�y��tvǂ�=P�1��7Rk����z��Ɍ�"���C�ߙ����c�L5����=��O�*��̸oxH)/�
E���q��<�;���A^wQ^V0g��R&��@s(:{20G�xj��o�����=��yn��"��jO�a-X}12Y��L�K�����	1���c�j0#<Ʀ�LD�Į&�_*Ě;�zll������=%��iMf�a����w�s�6q�.�\��ԟ'���efG�H_�H�㖢x;�ĵlJ����J녲QG���i�4o�y���5Vg���O!_�Q�3V��T{fx� ?�ß���5�P��o�E��U)����-w W1��J�ŲQs˗9�uTU&u��<�(��z�`���7l��O���d��Z�xb*۴�{�{�)\��)�'[;���:�aB�Ui>�t��;�m��T�Ho�@g����)��$�x��ґ�e�u�=�&�����s�';r��y�AD'`�<d���EJB�;f=�H(��b�����K�$�"��D����vN/��XY����׋��8��C�f�˽%�#'�5lҨ'�m<���l�o2.�`e)SX/��R|͏���x�;�"Tẋ���0�N���֭���:��zFq ��]G���������w�Z�Ok|��W���an71������o�{Ug��
�}9"���!%��c��y��MᎵ���}�<�̍��(�sk�/�iAyv�Z�u��G*I�d�	��r�8W�.Pg�6`s�'�����:E�k�-"�r�[ ���s�����X9�S�����8�=��@:]�'�ZI(.�Pj����~����GDѮ��䑢A�h��4������z���F_�~��g�dsE�0G0x^�s)\�4����E��ѝ�����Uy�<Kv���y�D̋x;�!7[�^P�#���	k�4�d}��[݋�0�W޴��v��l}�\y�!�zA��x2�6��ƺ��%v�Q:[�=~� ���j�����T��y��5��~S�X�#t�����Vm�����K�&����������j7hp�+n��g�<�@�&���C�o	"�a���9Q�*�&+��,��8)��~`_k_m�Ȱ�΢�S��+�J���3� 2��J�m���h�}K�b]�Se`#�����Y˵��[�y�����?I
�`x�d��SQ3N�F�A��|S����ى����m�Zz�'<���BT��9ۿ�kc��;�*K�F�H,6!���/���9("��21������
o��E�~�f[1i�En�����aCD�!A��B�P�(�QTooRD��lT�^�}�
�|y{t�)�^E��8ޗ�f�#3LsĎD�Q�ݎl=u�1�l�ma��0MvY�$2�h]�O��a���Ǻ;�W�#��/�P�%{�����f��D�o��t_ $E�ě��"�$�o�W����Z#wҬ� i[ɞ�[�C�F�bu!C�/� "/FV_�)���P�9���y�l#�6�B��]g�p)����C�Z�\I[*�Eb=��}�6G��D�#ߚe���w5>��"2]��;��8��n$mɍ�ȩ]��Y���`���Yj�k� �ʔ�m�-E��Z�E0�ғ"�=[�?t��NA������a��U鈺�l�t_��k%�X@4A������Q �B����y�֓�Eg�U��go�e�}��-�����`��t��(s6ID�PF�ې�<�E�Q% %oDJ�C�_��j��Wp_��@��4y!�I<�/�<�k�-8�ҟH�m��Qfs�^�lYD��7L��@��]���rY%p����M$���1�m�P���T�^FX/�2�E��K�*ԗ����G|��v���Ԋu΢6�R��D��v(���G��R��FR0�9�%f]��5�.���靹���e��C���O��
z�㤠l�x��Z�Q�Ke�AE
W᎑��+.#-r}�Ґs�{n��g�~��ђ���%㇯����ﹿ�\}h�w"�J��Պw�SG��������Ӹv/��j�<\��k�!1�='t�����2ǻx�<<���?��p�O�E���t�(��M��?�&��Y�MG��&ǎڎ�!&	������G��È�-+-�o��.�o��ָ�YYI�]�Y7R��MN�:�_�1�tD���I��<��l���7��z�U���r�i�#j�l�buQ��*a� lo�5r�iQ���:�`��*��2�ʾ{�f�_�M	�݉}�LZ9-�m_���F��W����#��r��~{�N?�5�>8H7�7W}N�u�ٲ����N��ŁX�j��E�����+���c�:���� ��w����<_X%�����/��X�������= �v����z�,�� ���-��EB�����b;�D<R�Q"����]���x�҆�MT8&dT����&w���J�����D� �pn����%
��1@GR޼\����hG.���V`o�8n7� 
��7@NK&�ũ�3C�;����A�]��\ތ��k#�6��p�C��)=�)���
;ĳ��@�b�b�J��]��x��w�t��O�#�b���h�*܃��0�a��M9���,��?���Oq��zѦh��zn6،W��G�D;u�'�X�v���唂zD>��?!��m<��ؾ�m�~�Gj�[��W�R_�<���$b��s �NdJm�s�����e�"�ђ�D�U����[�Y� 6d+��a?� 
9O)=���&�U˚�lݎ�uHhd�?���"��Ȓ��9~*�=�8�͑�&�����H	�ž�B�V�]��S���s�Q�[����2^�٣]�k�19}r�����:r(e�^�W3@��Yӌ�L��Gz���T7P���5x���[,�`U%��*�As�u.[�v�z�˗-��:�Z}*�$cq�i��o{����SK���T}�I�ۦ��C�T޸1�� D�l�U���n��*&�������S�ۢ*����7������h��W�����)���HJ��i�5
}pT-���e3ƶ��I6���kp��
�[���؍���JuTY�O���	�[�>^�n�@sZ�����?O9�$�]/cZ;b�<]h�l��!d4@��{�����2~چy��8�����nha��YI_�c���Rh)�|r��ܐ����#���R���$�G���`W�v�y��eH,��ڲe�u遃H���6�'�0���5�J��!�8C�.��
��lC�9�0�	�}-��d#�Eٚ
:�x��(�~���S�ҌH�^q��Ą���p��c�����@��*֢�_GM�6���K���W"M�B	_I�İ��
u����*4��
v���PPXg�H�L�j/#g�s�Z���wD��|}1�AK,F+�#�JjĢq�m��
�������m�OG �\��,��RЃ^
NƟfD�Wz��^x�z!�U��;���r~�=����t�qҎ\�������U���+m��v)RZ��f��@��_��L�.�[G�aǅ��8�E��xV�"�V��U�$�"ϼv���p��!�_�q��x'#��E����\f'�_y�Opp�v!Z�GF����\T��[��v��O�v,�M]��zq��7��]�S���x�o2��i5���~�]�v�,�q��=�\@���x��<_���N�A�����R����p߶Szj��U��]�\ND߻�O��˟�W$45�.\��]���~�Tg��$6��,'�G�I�r��L�c�ωA�9�:G�C� ���3M,�0ݩ5H�ޤ��U�w��uE��|��vz��P�<�o�c���Tl)�Q~�l���ކ{�K�P�A������̃G�v��U���Ux�i#�el�Y��RQ$�%n��x�3�<����Uu�Y���+\\��R�/�Q���@�K�{��zZA�o�ޮ��f��2 7�`T��U��0\;��
-$���TH���]0���4#��B���?� &Ըq��]Y� b�Ĉ=X@����{�
3�u��4<�5�d���U5��`O�F�,<,�kTCS2*�Yf��b{0&��M�^'��.�@dg�WŽ����I��u��3V���۪j���N%F6���iʟW&Y��#��ۛ���ɼ�G�%�$Fv/@��lG"����K�#�B�ݗX��&�n�\DT���|�^(���yQ�3��V3���PQu!x�?���f3�A�z�w�&Uڒf�aѣ�.�V����ƕ��r�{I�qj,��~(B���0�Ryܦ4!Ʃy=G"YUH�[uƉAo���*ũ�I<�T�_�rـ�[���]=�V��V�����#�Wo���ǽz,�+=y�]uI���4Y��ǹ��o�'�-�kqA�$S�s�u7���D��O�X�c�B���ϭs�ղ)M��~���QBl�OꟌE�fC���,�VzcF�^� T"��v 9G]�6�}@�gVD5��U�.�9}Ű�F�
Ծh.�;��r���u�8m(����z��Ge�|���\d�D��r�	gۣ6��Q�b���H�����"+k~_"�l��Ȗ�әTH�(�c]�������0���[�g�x`�k��)8\5��C�t��*����ߍZ���\T�N�#L��I�o"w 5��>�D��|mr�K�S�������-h"���(�>�i>�d1�!���]6r�+�
���c��l�J���t�B���OX%�!$k��s�?���=]v^��a�ݔ36���.tw� �DH�Q ��U����C uM1x&��
r�M�\K�yj��u�N�ٺ�*�HU�L����r�8Q���\���b�3�?�v]���2�^���Ħ֮�ф���I����ee��벳K�dP��B/�!?]��&o򅎒i1��!�":��-QfH�b�֘Dċ5��f�����ش���^�����k�"��3��T�d�����~��(�Niag��� ��V6F쪮<
o��ȡyaO��XD؀?�FfDv��SB}��nL��#���D�q>����Bn�l5e�¡�D�c�҈�0�Er� %�������+}���fL�[*ۦ�};�:1�EB{�#j�&��ʑv�w���g���x�׋rĭ6��]� ��uNG.Æ*}7A�����s��}�LX���$�£ŋ���}B+y�.-d��T~��F��:�e`;�mV-�a©�F�J$�[����uK����m'D�ݧ{�a̭ƥQ՛s�N;B�3��j����2>���1 �Ͻtq�|�X|w�㟛�xr�TY�������|%��P lC��.3)$����^��Nb~�<�=*id�i�nd��UeKx>ԹI�t�"ד�rh���M�Z�]U�����U0�p�/[U�a��~�*S�G��.A��.���K$�X�|gD����k�R�)�&O[|q�w�kb1�in�r<L&���8E��G4�VkJ�&�^c�����m#�2M�Ew
C�*��+ݕ\����D��]K榋$^-5M�1�=��#���a1Dҍo^�cX�-�Co�!j�s���规��Gx���lI����)k/S��� W��{�E�*��h��~Dlo:��(�"M��h�������
m�`�I��RE�b�UuP�o����0�i(6��#'��5d�I݀�s?��W{U� ,�VU�|@�*����+�]����S�,����r��\ :GŐ�x\�^C�$c��j����W*�6i4\��{�����|M~v�*�G6"�K��cYˤ�ċI~��k���rrE��)��i��|�ZB֘:#�"�H�zMӐd�=7]`�P��K���D3��SV���7�&��S6s�Z�KG��h+���|�w�����f)_�s������I�����&����<2����׺z����؁H�qC80;����rF��L(�݌�6��r�e��^�z>���w�J��9���
:��p���dFBt,d�1��1#��,��i�g��md=��n�.G�7�{*��_~n��ly��c�A�&��z�/z�q�ŉ���9C#��g8\�5m?^�Iq0JC:P�@�mg=�Ƞz�Y/�3(C���A���+S"Y(�%d,XT� ��@���m���@y�E�F@iTz-f��`P�l*�r,( ]`=���
f���[Y���_�px���۾��Ȗ���t�	�Y7�%p���_t|>ޡ�!q@b[ k6�E�i��}��X@�5yhdBgȊ��:�tt�����]��`lN���/�
$�@M��d���=���KGZ�[�tX*���~�ʑ2S멜��O"bA?1F��N0H�������L(�H`�,�L'�Y>�H�r��:z)��� ��9R�eS �2Ћ�P�N`�^�7�Z �Ӟ�`��Џ28��~�o����xM IsA�
���z@e�ס�^�@���FA�^���6J��X�!%���]����r[��7�!!$ƜaL6~n����4۱4�����.�jP�{u�w+L\���E�Xyy��Ɵ���WCUg�{%��Zx-�J+��ZBs�O8��.�i�����?�eLǧ%'�^��bT���1�y��mF�4���]pu���FX,�~d`[X��`�F�f�ʂ1�,�Øq��.�>�X�V�_�Lj��}irh��!��>9Q�S{D��1=&%)�,S:5�q�ʑ�	{�>��n�6 �,f�- +e�΂l��lBg���j�ME��/�ě� �8���H�T ��R0#)���p�Mt�Ft�7��m�IFtp�2�����8�-�����T|A��4ͽg|�e�:�B-�4����t<0��H��?���':V|kdv�?���J�t�q��`7c�:;듟���� �ۓF�s��a�ǣ�FR)���-�n��h22�ĸ��P�s�m;M������ �m|�E0'_u���;��\T<Lw�������`�DEL(��f^�c\m���+� ��Oǀ�Mz�Vu,C@�;O�p��M ���`r���
~+�$�-��Z:�Rn�k0��3:eB8P8w�NS�gƅs�н���J�]�LHt4I6.���ӝ�|���h(:��h-��e�J�ke�o�ŧ+��
ş��`�Q�vC��@rAрQ��5 ���v��g2�0�p�s�av*H���OK-���`�!��Kx�w_�孍��k8��-�5h�`�c����44�g$������-&3
�f ��e�{���k�����i3_f��з"�C�|8�����į4`+A��v,�8��3�b�q ��'�0Gf���eƁ�ǟ6�x�8��	ֶ`��_��-��>n_7j3t$ �m5F���r.���΂?~�5�j��O�r��q�QT�����Qmw��	& ����/��5�3!���#��	G�m��杦�F�ݗ@z��{��Go�K�L�H��K���ß�- I�	R�$cC^V�$Y���?rC������޽�d޸����po��?2�[����r����PK   u�XY�\HJ  �  /   images/57470e45-49b8-4c21-99d3-774ad112c262.jpg�wuTз���tw7")1CH#)�� ҍ
]�� �HIC	�)5t	Hw7<~w��޺޻�>���k����w����_ ����
  �x��9@( �������������������qe�c�gdd~�9������%����A =��br�b aBBBRRfrr1>N>���?·6 .�����$� �a<tk�>���	&�ѫI
�����������0L ���M�	���U����{p�(%�bb�oQ1�ejNk��I��c�J������G��l��%�����N�h��O!�ύ�I�$�xqc�>�c�� r��\y����u��l�t���9aP`5y�����m��x�������F��v����, ���%=Ӭ'i��=��ȿ��e2m����A#?LW��=}qd
L�p�yit��F~Jz�O�X����a��g|��� 1'Uz���v%/�:Xw�)��o=�Dsfw� cyf��r��j2�IA������v�}���+y�9��ԟ\4Q]*�}>w��B+w ��,���ߦ���V�vP��O
��;t�k��Ybѡ�Fw"H8�d���.��͈��2'a8:��P��G��c�[.�����,�.fhm;���ۏ�4�m�T� �S6j?-{�c�^��|�?v�O��O��݋ڸ�9z|S�C����a�lR%��o6VE�:���hg
ssx��"�����i����N���I3,�z�'����gbAwg��X�i�z^�h���	�2�X�Le/S�O6>[7ۭr�fp>���qx�ݝZ@����/�����l�ZC��&�%�8�|���6�;����2+�T����@�R��6~)kj�A�y�߅�J�|�=q$��m@p@�"yv(�O�}�6�*���������z�}߃��h*�
F�p�_|�J��#���Fѱu��<�FjL���i�7뗶10�p��S�o��S7�S��;�3�0lWս`�s�O!��K��ԉ:E ��/�W�ݙAD��<�A�x;%h^��a�&����Ζ�7@�xN�Ņ֚ИF��4f�J�iq�u��W��AA~D�c&k}ҜD��"�e��F�Rx���&���8�xC����֕� ٙR?ʭ����p�ѣ�=�:��Is?�� �La߭m��D�֬L-:Up���.�5���gm�M2t4u&<P�}���)�L����5"��0;��u*����:|8�����c�7��;���3Ɂܼ���ʿ���R�оc��!%/G���<9�FpI��2h<��dM�a�'��1�q�yC5��ZX����<�0.���^$ˇ
�hb���sX~�W9��ە�?�Gݢ��G��4m��>0P-.�G���&'�����bS�(n�ioh�&�M1��d�=7=�T��'h��OYT<Z��`'�«��b�6hU��TKKi�8o7_}�Sy ��M"�&Ŵ�"�M��Yy��8��G*1ʹ�ug8#����F�b��B$y�+N>2cL�c$�p*B�	���Fd$�n`ؿB4����i���f�n�җn��dEFH�J���x�����[o<�%5ba|8*�M&�����Z�A;���f6�a6���=�-id�����u���5?�EҠ������@a��w<='�뜭�z��Ic��1K�q.x�}��[�.v��;�h�/��}�����[ژ�%F�X�o���u��� �dO�q,t%!t�_���Yd��^�kf���|�7O�uvT�<bA	w??h��^�}i�?I.�M���=�����s˾L����ZŎ�O��0Hߏb��٨<��"����yb.-vAv�s?���b��ő0vO�� �=y��V�۹���A�B ǋ9r�{n�}�h�����M������Q�`.T�0�mȼa�M���@���j�*�AU����w�b��5U���ً��5$�����x���Z�Ǹ@���U���[��6�{sN9/>Y�U�`~z��?'g�_��!����
��r�" ���gE�K �a�C��ǲ$�s���|)�o�1X��&Qd.'~�yʺ���N���9�%����ƶ>����1�Is��WNؿ�7i�n:��R��y"E��	�8΍�}UTO~���8�X�'k.;X���E���2O	ʢ�)�?k���ڭ,ŋӠD_O��b���[�:�I+D���$7��CSh�s�#�J���K�7��ͽ�EF�Q�[�^XسTQ/� �T�u�;��PcA�Kjj~��05�G�^l<�O�^����6�&�{���>k��˦�L�U�V�����{�x��H'��X�,��\*ru��ֽ�Xt����+8��b��F�aB��*7�;��}@�OX�Da+�F�iq�^g�}��b�v0���s�c[�"\=�f��)S��";c
*��,�F�sR���26�����S=ް8y��֪�8k�����"i�0P:G�AUXON�I��#�-וTVxO���HԢU�H��1�W�V�K����M����,A�� �@�n�$��zF�p��ӓ����ȶ��M���TϹ��j��ͶP6@���;xE�U��G�Gz���*��ENt���b	��ߣ̈́���ys�.i5j�~�_?�c5���[UsK������4�e�1��>��6��)Y�<9q��׸�����k����4�W���+����<��������X0�_���R�͵pt�����5�澨w>���*Cahl��N�G}G��=��95�U�-�-p���C�A����hM��/�3ν�d�Ƙ�2ϼXk����>�b�2,�ӫ�aYuy>��6~�J���oB��4��;^"X�r�*k��Q���NM��c��7��$���%�@�w���L���U�ǇƠ��O�y�7a/�GL0~�8+�ͅ����KX����b��~~��� g
؏ԠL�Q3��{ok�/�_�3Q�Od�f��ٰ�!�ŗ���=���~ꂁ�c/�B�u�����6s�{v��3��$N�(w,�/y>��;��R6b���b,��xE�|����&b��A6�O���u����(�U4��� Z��i��NG ����Z�ٕ g���;׵��홫�xQ�<<�9���	:���\x��q��f!Тm*��S�8+b��3>Ea8��\�J�:i�D���#y�H����I�[��ى��Mv��$�Sr6Co��i�_��*j�$�k!e���;l\7���M�ۈw�
%vT�{(�� x���̆2��K)�Z� 2�Z����eG������sC��cg�
��f��Z���;�p��k�{�!Z�t}�Y�#r���gm����@��5n�a����D�?o��aM;����oS��[�� �ʋ�B��n���di�6s�I��G��p�21����J;�U�bss��W�k��n]�f�L����;x��MV�-���E~m��V�y���K��l[��1�$/_q'�}�&o���}�,If̹�d���-�w��f���h� �ԅ7�`����τ%
���3��e�8����?�hlA�K�˳s�af��g�h[Z�l�۩l~.���j$}�y\o#n�by�D�I���DFi�:6�#���(��>�����m�v*����B���8k21�Y��`��� ��ߔ��cLg�+_ן�6'�%EG�hX���e|������^���7	p8g�l>�{>��`���;��4Q���Dh����+@#�(.������xQ�H��y�b���=��E�Y����8YK�:u�_�uN�GSΐ�>�n��,�Ū�"�bA����p2�CKF`����Q�!��)�ԭ��uv!����Y�S��T,Hr���σ��x�ތ��4'����=m�+�L����U�r���Gt�S��r�[�������Љ�[�H�4���������49/�P��k4"��Έ�ȩ�U�7a��[� �b����7�wJ���?j�݁��1N�D�����^��u?��d��4M;�%>�3!�XZ���D5��U۝,�\����B ~'�B�E?�'aO>���׫��,'��YD�(�Fm:��'}V��˭IC1A�I�Ə��Q�&����T���`J�G�gk)��*G� ~�6ɒ�ʓF0yҼ��z�[�E���S��F)�?j�W:M��&11��;���$�XBW�g��U�O#D~k�n�-jx�3(�T9&���kP���3�k< �y�������)!� �\�����7��]K�t�d��;�5E�Cۑ(#��Y�����k�E�7�2�n� -�g�_@�G�Q���Զχ���*A�C ��u�P�ߐh�V�Ç.gpQ��f��֋�VX%�6��d��ʧ�	��4�����0�,�l@T�э�P�ڪ�RMI��G9I�ߥ%NI�\�<��[���OJ�h
g���L�a\��l�!ן��-�k��������e�j߭����A�S�I�6+dݯ��sS�Er���Lr�m�����y�l�x%0/ܒ_�Y��
�9k��c>1iH̓|�=
q-��,AxG.(����s����z=6,8�cO7�� 3��AJI�g�
}�!�]�[p�r'<�b�~���=��,;�o�7^��7��MU�M⣔J5��A�c3�N�To|/���j_���?� ���h�������˗���8��IN��qQK �KnM����b���Z_���7�qk��
��<s�x��X���'O�E\4<�*�u���U�^8�?��xS�M���(:���\�] �ۤ��(��B��.(<��^��\�{ H=r�N�l�e,}Ǌ��ص,�'#��s�+?�M��W^m�_hq�����q�}�H�_��KJb�oi��_v6!b9�!��&g�-��_��A�5b���_H@������5+SIAp�ʜ�j�(��W�$�D�yo+6L�=w�ղ�꾦/���썢Y�ȴ>�|'q��lk�FūﰻUT��a�u�Q�_;��`S�q�b~�]��/�	xM�#V��`.��w��rb#eg�%�;�9k�_k�}��3$ŃY�*tR:H����RF>/��k����s��<��J�T�'����c.��Ң�pV.���d���������c�ڿ�}RF)h�u���޹a����:Q����rh�{v��2��� ��1�<�V���ʶ
�Y�~հ������*0�f�����"�rH�2;v�>zi�㤦�+R�)���y� ���nJl�x�a�>��C��N��~�n��O:[v��)l���ę|oX��*
��mMA��/CО	����e��t�:����̄T#+y+2G?���е���l�gr?�����w��Zas*A�⼏3p�Q:Oj�^Z��]�kd@��(koo�㧌�o�#�Eg��-<Z,��$v��!mM�eą��>t�p�ri Q�6_[�����wx��_8�?��&e�3X|�~-1����_�;�9!d9;�x 4$�T�D��E^�[����Z�B�^HF(����c�:Z~a�9۔B��^3� ��G��Զ����;�[ͅ�٨4q'o�K��i �����eSHQ��윻�Oh���h�C�)�}ŕ􋣕U4�3(� ���\9���у����T|"#z�;�e>o�+�ZG>]�*�?�Z�V�A6<��K?X
Z�Z˚�H2� �i	t}c����=����paj��Α�)�,0_�R��W/������mǪ��k%�ʎ�7:O`�G#��σ{j�X�ǁ<Z z�R%KQ��_G��ᮢ�⃍w\�ĹS2LJuw5_z�����u�=C�ޱ \� �c�s�s��/	Sz�0�țwB���l_<)��T�M���݋�n�V;]bg��N� ��7R�$��`�!_�9� �S��!|s�#ςԔo�A}P� �i`:p����Wы�\�AOOv��hd�bQ-P-rO��0�3I��8�7"�?D�$$�||ebzH4�ς����)�>�!0�$�3���*�W-����W�h_��6<Q?�.why�[����rt�[�>dYQ�&RGGL-U>�lټӳN���4�4;��1?g
�����7�Dq,4T ��gUm�ܤ�j�3������ |�y�&|I��`�uEmQ��#�s}� I��=����U�� e�e�Gg��,�g�$Ei����$�6�[c�s���T�B]t�)FF��}�}� �0Y��9!Y<VV۾���5�28�3���62����yo
T~�r�B��Ab�)���o���G�v_���+%5F�pV�'ʵ����_pU�T��;��P�.4�v3�����,�N����"�)�Yn��P=J�6(�~7G��x�쨣��"����n��R�p`�b�۴�%&�n�5B��8��*ɒH��|T��j�X=�U$�c����$�Z̀Г�&J:p� F�A�������[�_�J�6���b~:�a�^�89��>ў��Kݜ�[�AŠjqߓ�f�Չ�<��$���.���<��SUyI�2�awQ��t�$M��H��P���z'\�M`��6��@��D�/��}7x��f���H�4�/y"|,[�� K�)O[pH_��s6�X�5�D���	*� ��6�Y��4D�h*�����7�M���3��$3�PK   D�X�Rr5�  5 /   images/5dbae223-cfe3-43b3-aef6-7502dc6b2367.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   D�X�@M��  2�  /   images/5f70de14-173d-45a7-8b46-cd4e4e8c904e.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   .{�X��p� �� /   images/7e81f6ad-0912-4ff6-bfc6-e58bb7840941.png�wT���6�qPDG����>� J�@��R�FjpP�A@����& ��&���"=@BB�{��=��������z�g�������>{_��{�s􅞎������@ �ݾ��>���`�t�����1"���mã�8z�9���>�e�@�|�9T��� ����������B��=tu�yd���!��p�8��������_���/"_�c�?Ə�c�?Ə�c�?Ə�c�?���#x��ap3 q�1tS����1~����1~����1~����1~��+���������f~��ռ�䣊ʷ���������N��W�e9��;��Z�����=�����/�̍.����;��'��Xb������jR��Rӭ7�_��tg�WQ��;G�v77�Ҩ#�S�v�P��d�^uw���wE~����1~����1�?��C�qLw��J/i`���[1U��*����hqE��R)Va��jt˗/�,vLe����|�)��*�N}_CW~�����C6om�Iu��Fo]���O���j����Ӄ�adF�� ɜ�)jϣ]�x�A+�n�iz�����T�'3�Ԑ\�c�t5��^�ih�_͔;�o`��&����Y�O������HA2������h�bw�χ��k�N�>aS�淟�~B�Du����X�<�a+l#Z�V��yf�._{|og#����n��Q����:Í[�(1�u����I���7�<�Η}繻���_��ƿ�lB��Qx�ING�^�Q:�`ݦfB���úL�?b>߉g
gVO���$���d�W5�p��s=�[�-��d�z%��`�zd�����S�
�2NU���go���3~ϋ=��#��y�-�-� ߹.�2[��.�u,goz�&
rZ�T��88���<��Z#h_���İ���uX/�sTF�lG�h�[��t�ڈ�i<��3\����e��o0��p{�R���O|��b����t�� Tw���|�e� �')�^��1�"�c�Y<�-a3�ç�fV��A�E@Z^�S^�Aś����-�_�b���a�C�䩡���&�@S=��R`�/n7u*�K�f2����z�̂*UR�Xw����;J���mIW������Nz��p�l�;TmV��Hi��&f�ee�RX�_צx[��6&��4�7k=�k
�P��ah�c�{�h��rvv�����ͩV�K�Ֆ1;W�g���s:�8=oQ>~ؽ�|��["y�8�d��9V���m�T�Y҂�_C0߮mH$�;.J��s'����X�Էe�:Nڥ��R1�?�dV���+'����pזA�G=���3��NP�jc:�����f,� ȳg:<k�\Vj���U�b��h�zE���n�(Ѱ?%eHm$��:i��QyuYK�������hs[�9�v�E�}#��=AYɚͷ�����j6��~����×�j9������%�I�±��Ð�m_X3��٥x�6�4�� �1}*u�:6[ĺ|�i�CI�{K�\��-�ӰO�� }�/}D���d1�6�Ű�Z[��
�}G�2OUg�@�\��n䊳IKA����	��~y��]��>��\7�(�qj�?ޛ&YX���Yf��קּw�r�e*�)��Z��(
|�KI<񓳨�r@]u��5o��
vL_d<�dL�U�և��R����T��@���_��}橒�b::c'h�m%`��t#߿��B2"�'�%��+'���g�ZT�+\�y"j����կ^�ʙ�P����#��{�ld�p1�y�?3��˫.���^+�Zm���u`�a�Z�]��-��]��PA�9�}�z��k��o��ru����i�&=����/(��}���!O�Z	�gg��oQ�7�	�������n#�~1��|ʘ����~7�����V���Ɗ��<yD^��bd=d'�S�$�^L{�ؖ'��1I�v��˯��uYW���Gf�U0"�뱱�u�2�ל�����5��
����j%�7TKj����6+k#��'��{L[~�l�5��	��I��gU;u�,��r�{ ~ G]��$+(Ĕ1�VQW瘋�r5sp�tv�:���n��������%����0�)w9ח�rRRO'�\�|Z�A Ѷ���S1�ڔ��	�@�־Ɉ\]�tV���6��U>�WxG��n�>D�J�9�ݯ &UlX�Ƒd�p�v�a;Vb|�l9aX?,�y =�9\��yI�/��|���Y{ٹK�"��Dٲd>e��k=M2(�R)	�t����A��|��A��msKd�zr�V�@Gk�
�ѐb��m{:q"��s��C�SY�n�U��`aف1ȇ<����Te?K��M�;��Z:�^&��G�/mΑ�s�ܻV�h��{x�}���;�Z�B�~K��ʻ��	)i�������d���:o�~6������s���
���((P�n���ӂ�ac���l`>{�8R��l���+buڶ�j�V�4���9�,�ys�ҋ �R�ᇠQ�.��m��~���ѥ�KYLO �E�<ǧ�RjG��د�_iV���:F��u�[mqkG��N��y�ٷ���	���>~�b�IDW%�*a�$�]<�Iſ"�D\��5m��F̺���n�u�S�I�,�c�U�B?iɇ�	_�'Xơ�O�8Bmx�̧�u�֫��<e[�\��b���|���{�}���>�Xn���E;�Z9&�,͉Ц��]�m�������a�7�خ	�l�"�u��YsHQ'�{g��=��ItouRz��ϝ>��1Tc?d]���zJ�LE�C�}p���X�1�I��.I�J��55Ͱ�lw0�X�Ī��n(RSC��=Y;��ۙ�S�A�C'V��Hl;u�PT%v��١E+X�6�F�H vt���h�I�M\I�&!��/4]ޚ#w��.+2h�(����CV�.�8����s'�k�IY����� `�b�K�)V���UϧJ��_��x �=h�c��&BOqw¶�w��
_!ƨ\����i�X�>�ғ�+�u�׊�wO�y��S~�B��ߦy�9�yI�.�*� ~�x[�(M�����3�����ÿ�󒵔(s���my>��7�C��� vx����բH@ɋ�Q�w�)� ��A��}�Fw�b�+����U�^`au����9GR򘲴K���ŊJ��n��.x6j�����j�s+�g�So\��e��Y�3~S���1+$��j]�����&{hnTM��=��B幖ۗ�k� ���џ=�+�26����2�.�
;�d�S��(a����3���#:�;�K�wJ���Lŕ���Z(�w��Xѕ��a`ZBy&8�v/zB�j��"�i�ig�� �����.��w�eZ33�)hb��< QIi�P49�]<Cq�,��,���x��@�>qJ1�g/�,��zѿ��@奧P�N��*�_Э���ج{m��:H&T�����I2�߾�S=a.�p�tX���S}�]d|�д��P�su�Ǝ?���*({&�w���l�ZHClP��1�S�tMzlMdi6���k��3>��T��Qo�^�D�1��ޠ�~K��]V�w!ҖK�j-ۃ��Ui�뽷��W��_���X�9��0w_��Si���.�s`��Dn]����y�7]̑	��E����
U��>@��9|��7�	��k��s�u����RJ�3> I9;��nށ��0%Y��卤)u���Q]�ޖ�eđ�߳|���bg+��v�O�欪��9�2�� 8��f6!i��}�	���~���VC5U�0T�����+�*t���@�K:xM�bt��ux�lܗ�&BX�ˡ�i�������Hߩ�#�0�FE@vt�:c�dlz��$c�k��2����0��B�m[��:Qy�Hb���V�$�оN��jc�_�0��CB(;~Y�4@��^��ި����>%�S����s��2�ǯ�D!vv��ؐ�1Z^*�!���]�o���z.������M�f>��琾�`x6���o1&�-�;|����?o8r��x2<�c�Y>�9��a��q��T�O�jX������38-�tN�~5M����2O�}�ub��ޖ�0+�����m�uv�l���1��]sT���APH�� d3�D�dQ��^��%g�>e�x"�)�r�b�H�
Y#�"iqYvu��|�����FZ�U\�!=�/`F<��v57/��2�g]��������z��+��&].�p�4e>\�L��`y7��[�!$�,f�k�}=�Ņd=HM9�F��+6��hU��T���A���+���..�����Ld�CjJ����m��Qƿd��2��avj���t|��������XGd��"�[�FN����ؼF6����@�g8$�)��2�����fKU���A�)��q�����$��,�iO@��]��L�\>k�V�Q_t���6d��F~�O��S9�K���& �AR˃�"��S����1�!��S+
v��������6��23|�{Qt�!E�eN������
�{�� �dJ+pȼ
ӛ�������3(?�V^c��s�����n��B`�u��7~S%�Kا�A�+����pp�~[���ԶV�9�~-���
���t�2	��VX�g(�R�M"�?�	@�uGJwK��O��X��YڭU�C �VС0lȖ�B��V�N�f���5�����N�Eë�﯌����������$Ɲ�����
.����^�ŏ�{���I��״e_L���;����Q,�,����8���!��Rkq����Ҫ����m�r���]i/�?C� ���"�x�
�8:ٰ!�!��r� ��_̻��ϊ�cx��)�X���D)�� s�4�X����}�Av��,з��"�7��{�P�oU&�o� ��RQ���|e��\Eo�N#2ԑt��/fӟSJЯb{�¤,�C9p���A|ښ�Q�.U@�;��>�ttl�V"�#6�!%.8-V��@��@��W�����E�V�UM%�Hn3,/=.t�!�����!P��W)C��֍�,p0�b.#��U�l�Ыk}mTz�87�6!�������W���F��BWͅ�r�4��[��Z�sdF�V���IB?�c��`��/��1,WD��')�o���x��7��J�6�;�n%��������!c�5�\�ñ���}<�W�yI"�*B��}����,pl��Ímd�C�S�컶H��z��tG���\��T{`a����ۈ�Pes�i]fS�;Yp���-�/�/~�V��!0Rj�=]P��ҏ�=�|���+B�#��6�s���������/�aH�'ݴ3��@'O	1�\_WV��Em���0�����<���òx6����U��l.���&@�,<�a���=\�Ɇ�	�W�h�&s�@�ջG�#�yow%rE�	']1������E���^q�O	�r-\�;�?��4�� �'��>	F1� �ʓ����jf�9�Ĉ�&G@�Gj��KY��tub��J�N&.��#B��Y��铥fÉ�Tܕ7%Ѡ~ַ�r�9w{�7:�=��Da�WC����[vh۩*�����=����l��V���LʴC-M���xQ�Vj�}M�<�&�C��}�='�KB���q�5[je"F��T=1�ҥ$A��D�߆�6@A1������F�{%2���3j�u�E�Zˊ7��2*�g�v;)_��i�rR�R���R��/�]n=�C+ԖWynU��Q��H����>�=�S)(�ڏ��r������I,���&�(ut������I���q<�Pr�*ЭY�մm?��t�����&�߻�E<j�/�8�o s@[�_D���Ed�����)9\�B?D��V�G�����YU��������%�{�-�R���&��A^�"�-�����X�����5�L0���/@Wh�����T�c�mϰ�+4#�U�����x�`�+���6zH��yaڃ�ZL��%o�<G�;]�?Qam�vg9)�̩��΢�r3��؏0x^���'`�2t���.� �*э�qz^:K,��T�z��	R^��{��oE��}R)eʎ���lL�Z��}��Z�Av�m��^z�,hH�w�]~jv�n��7�TTu㴙�֍5����?�:@&k
$*�#`K[�E�]����H(��@#�J�b#JDNя��8oI���2Y5q�!I�w-�ha�ns�2`N��������Kc2%�p�=Z;��R�\/%E���F��G8�&<'5_�%�ғ1�u76e�� d�!�	3��ų���"Z��X2��`�wfIW� 
Yv�,�
�^���b��X�%-Eos�U�ӹ�vބ��I�A����c Z�?��/��R�7Ǩ���]u����G;J\"�q��_���zǥ����t�2�M�����j�hw�Z��"W%�j�d�L�)��q#�*���gA[��J&ٜ���J�6�W�d@�g'|ͮH�\�{BnC9	��_.�,6�^;��?��Y(	����+U���ŻX{�=ڐq��.�䲷�x.�k�JGb� ���rK�A7ܥ��}�+�� ����#2��������Ak�vf[$q9%�<A�b\:�"<e5���J�������$�(��B�X��Z�JĖ49� �ڃ8�!O��ϵ�&FIb0�-���[�<��n�U�)����y�y"������l[KNEgF>���@t��eT��0n~�����Ģ�zg`KE�@�� ����z�l��o/���=:���4?��Q��st;����m_t���n�/�yP�2���/�o]+�dg�\��X��;�>��$�,��$q9�f�ʩ�R�oA��>�����}�Cg3�0k4r;W���W�T�<!` �r;hv������SP�́p���:��Hն���H�Qg��0���M +n��4w���E>����~i)�(l���T����ڻ�q�M��<����oOOeAC�W��f�)j.Y���b�{��y����<7��6.Wák]b>����of��)����Fa�Q�qګo^�T�JӁ�A�'NT�&���T�"O/hᜧJ��襕���y
B�Z�:$�\F�s�7L�&lϋg�󅹦�؀�v'Tv'��ن��a�@�$���q#S|üDx	R�z�Hp�ޅ`%�?q��_,�!����F|�*�����9F0Mw����u�u�w�Ƶ>��	l���D����}�e�n;�I�*������?IN59`R'(QE�����5J�<۪�^����DHJKF�v�[S}o�t`�#��|,7��k.S!�A�$�u����E�|E�Uȶo �b�26/u�
�[�P�tu��]} �3��;�	�}������+��q�eؼ����������9`K�H�99	BQ�a����rZ��E�FN�US'�)�t�s��GYHZ��j�@Ep8�m�n�{���C~�ӭ6�~C�v�I���T�
3)�4��s��%����[���^� i=lS�9��S�
���o�װ�@���X���Mf�Ʀ��O�����[w�N�v|�ڊj���#8�d�!k%$a}�6�;�i�,i�!C֭���X���� {�Ta��7˾�$?����W�R��AΕ���ef���H`06C��>�bn�"�<q�%�1�p�bDX�\�Ɏ��8���W�P��<�|�/�Z7���ą �����>��}��4��!����P������o��	F��Mw��uu��X,�88�5�i޾�cfIs�"-x@`07�T��Z�G�� �#���~�m_��T^b���Rg��_Cs��m�A�f(��继G�*Ქ��{�w~� k���M�̆ {D�KY��+�L����'9Ze%�#�ۯ������%֞��|�4IH�G�@��y~\⎛4����mp�r&vGƫ!,���"^r�
�f�դ����Y���(M(&Vo�ncL�Ғ�~i}�Т�*�ۃ�J3rW�P�+���\�����|v)pU�r�"��s����7m�w�H��y�<�Nvn.���*�;���y5W+�e�x:4KH胝�p��8.b�����jJ�s1�JNn�	��~r#x���_��Ax	�o��[�$���b�nDM֢��9�%��3[AU6l|�B�{�}T��Tx)�N�*�@\s��U`~���a �����I׈�h���c�0�YS��o~������?��|J�����^�n��T@��ϪO�
4���g���|�~ڢ��q���@^]�!�P���`+R:e�K!�?�5���E��xuQ� ��*�!��] (pi�t,�֤�4& ��zk��]Bw�R2���X�c��jlbo�ѿ˿�r����SDt�il��Y�t�N+��59e0�1^;��}>\J#O���p�a�Uk����CV�G��ҊP�:K/��e����P+�*ׄ������ֲ^�aֺ�7�6�GŌab�0Ъ�̽�>��2�	����z�+\'.���Ź,A���IaR�G(X|�2(��٫�������7�r�K��6�-��갲m}�c�g��oħ��A�Z��ՂD��^��j�`#ζ F~�_��b�@��k�	���~Nש���Pi��8�+��ey����@�.��0V޵�oJĥ����� 2�c���	4�E�����Qq�SdQHOF����r����T!��9ed�`��4��,�BS9X(�۲�Ŧ�^��Mr�8��{.�\3�š�M��=Q�[����ZCZ.|r�-�=�3a�+�
$���$�g���B��Z�x�@��y����<k͙/|ỿ�����W>��"/�u:W=K@��Hm�8��e��x�U�-lL�LL�KU�0�I�,Ts ʛ���)�����_�X��=n���`E������s����������s7��K �Lov�����J���e�M,�{�in���}?*�/]=�T����������G�'_&�m������.Bg�,ъd�+�Rj.���}��M��.ּ����89�a��;ݩ�*N�ʝ+W[w�n�Y���� �M�h�tm� ��5A*6J��i�m�O���3R9kf��b?-��N��b�{E���N^l���U��>��*y�;�y:��j1��'zD�2̖�� S#�F+]�D���o�bw�֬��Y���K�F�ϙQZ��Ҫ�,�0╶K]��Ֆ��EK;��M)W�%�+��NG�i���Ҍj�����]�@�.�V)z�G��N����S6A��ז���B�@v��s����\�W���5t���|���Q܉�;u$�`��"۫�S��I`�+����愰]w��/�u�N$����]�C0�L������i�~�Etb����0�_��5đ�����6SS'ǩ[m;a���&�VO��]��(�啣5U�<�z��O�F �Z�;���5H����}��c&�(�7K�Dy�Q��A����|Y�?M�h�]��]�aT���.k@tQ7�Hս���!��hڙJ@��tMyj�~���� ���{^U�4`}F]M��Җ8q!a����]<h����.]�}]�q���G �ܑy��c��2���&Z����!�!;OB�M��rMR8��|@6/H1��&�ϐ��_���=x7f^�w�11������ܓ���8���ɯ�5���-�n\��R`"�a��6��X����xJ��A��J���J��e&G3�/ӆbё(q�Ͷ�_�8��i�S��Z�b�:Ӭ>�ޜ�B,_ﾶ�GIϗf�\W7��MV/]k�G}xh'����!�"U{�s�Gną!%�w�M�A"����B����\��#��Νl�R;��ouGSӦ�ŕ�İ*�GP�-���D#.�nD9N��}L�@�:����<|?���ӗ_�f��P���G~���K)�?צ�Jg����&��Y+�	�#b�7O�[��u��an/�
.H /�bx�U3�C���Ԑ�\�eC���ʉ ~mJyx���X��_��
(����s����p��l�蟇�s߇��c�C�KAx���-�x֓�#o��p(瘁Zr��>�B�F��r�������)�����0���<H��1� 7��� K0�Y?�iV�&�4�n��o`1�$îg���)����#5���?OX�xdd�&͗���w�Č���A�g욍��|I���ׄ��e7&�#���+~�$D�cު�W�C�]�5�۝ SZ���`�۱�"V����␙�F��(����ް��qbזW��vg��)*EFY�?!�:�Zq����\�V��1�|��B�E%���ڝOimq����?�w�]�UA�Zrm���@ċ���!�-��<���3ޡ�� w���'B]ggW���:�3��Q�Mz>1\9�GT*�P���+�S%}�d%R���^�N���8~
n���UO2�۲bo����;��C��{����O�YM斏�,�½�)H�b���\�X�mZv���q����o���M���t�ҚI����逘�炦w����&�\j}��`"ɍi�r1�>}B�� ��Sw{K�9>��sb�It��?J�Y�cvs���q�XJ�iS�:�^mЀ��>,����{�zH��Eo&�,Ɂ(y1������2|n�f`���1��������O�­v�,ب*�0�I5.�=	n0���8D1���)��.��V�\�ͱ�����U�B�N(����Ş�� �P�����}|�}�Aum܄��%j68��ً5�����1�v(�w��5�3A.P��'/\`��^A�s.e���A�V�zG������j�zt|�����H�]�c�F����ۥd�T�-�:��f�*Պ��ֱ>�yϕ_��ؓi��MQE٤I1by��'ZDk��y��i�%��k�0�C}�?�gA�{�����E9,�~v�<cV����ͭ�,��Iхvvw�"�c�����Xa���t�ڶ��7�[B�h�@�Ã��#�$����L�U��b�q������!���G�*�w�-���y���^���`�څ�����~2��u$���>�T	�ڧ{��>s�'|�b��
ǑMZ��d�R}�Ě�10z��y�>״������4z_��|![h�"�=��:�J����I����ڿ��6��X���Z��������]_�ɽ�g2�Vh�+ʑ�%���]P-���4�6��-8��Gd��s����M\�N��(koG���$���jCdM���V�ϡ\e�GG����_0��l.8�~����<�$H$4�V�N�b읬��&���ʹ,Ƕ)N�88/�������Z��ú7_����}���d?R���T��N�ԉ���b���'�>�w��ݔƒ� vV(߷90J����/�$l�(u������꧛����IO,��&�Ʉ�/�琿���\��(s�Q�RN�ء�y�����l8���o#���<���P�P��>Kު�N�lDy��ҵR?�h���n�
Bkpk��~��L���TT�{�ې�ג���{FT>���M�(�t-��#��sȪR�����x'.�.,*��|h�z����eܾq8K�+7�p?�h�`F��N*`��By����Den%Zh��,�
|�����V����Y=z����#*d�,/�����M2(�	�g�I"�M��C����%���wA4����d��#(�ѷ�m��/Ʋ���6��#�����Ru��Ø��e\/3�K%�����C��5v�a�{�f���qU�L�Q��LC�^����G1f�A�jʡ����qyLz9�`�:���oC���np�����[4��-�SmzPHW9���l�32s�.kԠ�2�n	�)W�u�cu��&s��k����1�l�P`ey܃"��ࣽ�wBM��`��Y6ʔ�7S�-�AhӘJP��r�5��G�\�	0�eAZ@β�>oo;��2JƔ p�]�I~���RQ$��'f׽�*7�\tT������i+W����%s�`� ﻍ�;Q:�]�]x��K���M��&W?5*T4o�N�4 ��\�Bp�z���] ��H�j�gMhg�B���W��M����,;x5�cU��okx���(giP�+*\qb)���P�49�qpn}꘹���
� ����)�(��xZe�%D��u���Fe�KF�ċ� �������O�%�BY���w����x��cP�Ń��A�Yim��h3H����|}7�Os杖�ݤc��ς��LylM�w���D�KE��h��b��/[8�t���<�`i�����Ci��jx���2�֯�Gy�^�J¸-�KB��U3����'��*�A=r�<j�s�Egכ*!�l�3h�6rZ�������3��K� ����Aש(&���:��y gT9�X���/
�	g�Wb�k�~-��y��=�7>��JYҤad�� D
!��',��f,Ɂ�Jm�rv\���a]O��;X�0����Ѻ�l�L��X�A���b���3US,<y[�=�������=gq����D���ej��Yo���Pҟ?�>O�"eD�MP������&�x!U�̂���S<���5���]�	��>`���KobP>����Ú��Q���RT���@���<��sSy/A�O�,��X�p?�a(��x\�9οv�W���sH}�i|���U��
�@Xx<�S�5��1oTo<m�A�Z�����T�X}�լ'ʝ���--��?��O&6�f����!�M>�"��Y�]/��j�q;�d�Zl�����[���[[���Q)�In����~7�%JJ��kr���yd��mȽV&���Th���}�������R��"������t+��t�r���ky)��F}#S��H�9�2�k�\�g.C'x��B9�ذ�L</٣(�q����>w'}	��;|d+A[�o1vdt�y�ߡ�i��a��By,�`AnfJ���;>5h�^�6���ŭ�7k�P�;���*���Pe.��8H��6I��xm�#��������CQ܀@6z(8�m�3i���s)��T%�W���ߦ,o;�&�9,�
��%���>?��
���$�@�y٬�r{Kß��i����U�����Շ�^��?/U 7�E�99�n���}��|	'�z�����dP|�PG�A�?їȊ�%�]h��tMv�{�<U����
T��g��U�)�C8��I�N�
 �6��e�s!��j#c�6h��h����C�C~*2f/+�D,�3����{p�ǃ�		�����������\39�?��ֽ���5lФ�p���ŧ�y�Mx����b�f-�=�[��v��PlH ����~�_�R�';k�R>'+��T�K�>'#l�6���!0�oBm�p�g?̕���Ĩ���Q�1�ʿߌ*�$�;���/8��Vb��~AN�RZ��6�DU����c���rS��i��rF���{ْev��Z�Cm�x�e�d�Jiy�- @־��c
߿�h�վ� t�g0�\ꩦ|�45�o^��1��l��I��qe@���ݛXN�j@E^"�v\��������ֿ ��7Q�[g���{Bi+_��R^�VҴX�B[h�!;(iZX��Y�Fz �+��JH���PNgK��*�F{�KI�.�oC�.�`)*�"�θb;�v���\��f-.����ޓ�ҡM��!���e��P�"neW�d� .��x�S���^�LB�ƛm`�L%{��rVf�.�s#e��y�]8��w������2��6�� ��{�$N;� ��?Շ��-�^��Y�py\�ɺƦo��d�]6���x\���(�ȟ6��^H�x:���Glk��������	�]?�&�*ja�D����p��RO�Z��v�&�u(�L%x��&��U
��ѣ��L2�|E��oweZ�����Q��i�i ��+�J
Wy�tH2���NW�er����V�ߟ����/x�V�g4j���˳c���;�`�	��}g���n���!cpʖ����+N"Y�q�p(R�nP������k���X���)��Π.���َ�̈��ܰ��NĚ~�4'�,P�(����03�����n^*=Q9����m����y�RXj�s����I����&*hO}�g �Gn̾ў�_��
��U'��c�Υؓ��Ը�eP�
��G�Oơ��^�ল1d��	@�ɻ���YY�e��jԊ)=�x�ڷ��xx�	^n9�恃U�'��w�	�F2�-�%܍x�=�I� ���Xl���V F[6�����b����yo������n;As��~�-��!�%y.QcV@�G3����Bӌ�񔦇>a)���y�9D;P@2F9�<C�#.2��q�c-N����w��h]��8�����`mNy��:��������Mى�g�I?�f���GS)��ON>��`1WN�('������d���ۂ�L�x��K�"���Z��3C]�g�:�GD��� KP8�ɻ�!�85���ʁ�\ t��e!ȥF����H}�}|侽H��*�`�����<æ�h���P�~�c��	��A������L�YY��g���*yk��^@���TV�l��%Iy+%�>�#��1w�_O([<��[��标P�\{��=3�,Y�#0MҔk�o�\��t�*�d�Fz,e7}3Zڥ��|g)pe�!�n�������垠2�U�sb��%��
���3�'�3d�/�pn�x�����"n:`kt��ʃD�Lpֵ�>�j�����Ã�&o�GS����݅��ӛ�7W�6�=m~�A�W�K矉.�51�-��yzB�-s��������"�������"#��4��ND�A'5�����O�uC:�� �X^�%١�����'TA���Pn����KOe��cN����{�6�#�bZZ���x�OvX��|�/���F�*����df1 �V��*�R�~���׹~���q�Q�{P���fȐ[���E�Y��$��ģ�̨���Q`�\����g�Q>/7���Ɛ�Y�2���
�@��$��kt'��S���	��6Zw�e]��bHBRD��~z��NHbe8�({�BPH}�^#����+s����yx^�l�U�L���^���%�+��b�a1� �����(���E�R�H�/�|�/��u�)���y=���_�t3/�'�Z~oCzȏ�O�|�i��#��7�H�F����.�&�_oOA(��vf�"�lַ(Qp��?�y��G��Q����%�oP"~%r���K�!=vÚ�����v}�@�y�޻|�����3TK9�dχ���F_�bT���b-0���=��I�zK٧�1V��u`�$J,d�q��Ժ[Yf���5,Yy��-���L�`C��^3�ڍ
<D�۠���,v������t�|�Ir�#��!�X����7�bF^R�@�����#G]ï�2��̯�lsQZ{�'a����7��M�G'�cR�:	��Sߪh�׎�*n:D�~�+֭�N��>��NL�ƀW�8�����bl���_�>�8R���=��v�s�i*z�P�I�0!��I�l^nU��%��/@�fFa��M-MWK�Q7 Ӱ�S��3L�'֨� ���f��kD��i�͆��1�b�D�Ƿ���bǔ�
�_v���DZ�?�G�|g����ݏ5h�OL^�l�?�Ht<��x�8�d�����>��/_k!�
GH��{�9�������Y�VP.�/[���3��Zu@�rƎ l�v|P�`S{I��b�8di��g��'m��j�.f��}Q���F7�~uD �V�`��4�x%�7r�:�)�#�C�F�����fW֧$Sp�,�!8�7�(BqK���^���^/Pכ{vI�p����x�X
|}^�K�7|Y�׫�A|W|�P�Y�t=�L���ʗ��<�fe�+찳�p _�/rlr%�{���������6Kl��ޣ��8�8i�c����I��c��g�3��|�]Hŉ���i�i#&�)x�Z��
aݸ�z��ґ�4�4�n���z3���K#+���=[xf�<�"n(Oqs�k��M��� ->�U�f�~;��y�%h }'_��p�T9�2���c��$����x�&޵0Ļ�g�FJ=��L�|�x%v�����	��_B�'3�����qd�ЫU��'�	��>#�)�̛4͎�%K^�Uff���6O�^Ȍbll��Vs��CUF�X�s�i0��1��W*Qf|ڟ��A`ˋ7WLa�����r��kq� ����\��͊"�3$DS�ޚ�7��+�$0��)Ox�g�Q�AJ�SG�=��{�U��������o�Y���}Ė'�֋\<E��6����n��-?n���5i_D�˒G���E�P�&��&M�/��Fs��{kS�ʖG	 ̾ߎh��G�ZR���-���/���ٮ�f�:� ��=$}E�$:7��T�i%fJ
�/t�'���	ZY�������po�+/��_�r���=�a3<�
1њD������g�v�7��>(�0!/�_���)�-�B5���:&D����#O��am�nE!Ȣv��w��O�]m��S����Yk�M�'t�E\�<H2�`ȕx?9�@!Ӭ9�PP��n���v�y8 ��_rVZ)�!��Wd)�?x�nOH�Xͫ=">]ʊ��\�s�Pv���p/.��j�3�(\���6w��]��/2�%����>	��d�8��R��5>�����6n�C�#%P����o�9Q���C�~~姧�u�]�sN�"�o0!^ł���ӁSfeߚ��a�3�sn�a�9g�2�[�VX*��Ar°�V ���*A��] �J�fOH��ߛR�2\
um��},���8ǎ$_�l�y�=)[�dN8!��<@��@t� Y�5)���x����q�޽�5K\M2ȧg*�H�&s�v��_s�����P��FX�#�[U�m:�@%!���HVOiDޭ�S��<�e������u�s����x�?/�PI�xl��� ��T3�=w���7Bm�v:�����K,�ryW �S��v& z��%fY��rU�i͌���&8Y��۶@Ia��!][�,�5����$��z��I���K�'�-�3l���:BCN�"�O�6=�m����ό#�����{�E~���L �ĜV�X��u�uK�Ce���� V�|���J�)�/����U�����m�x[�}�ok�=W>�L[*�����k��4�4������|M!vC"3���_GWW��Sރ�<P�q����-g.L~��*a�jB�}�Gc*�����_����0��:���2Y*i��u�~<=�^°��C_���Ղ�Z"΂
|�������˹@��>1��A�2ű�YI�[j�eJ����Y"�~��!��� Q��=x[������D��D�\Hݔ�6�#�R"��c�����R�瞧	_�l����J�� ���%;{M�ه�+FeQ��(�b��Eňu��V� �M��4�8P��:՝$r���c ������C��o��8_�X�(�Z�������LC���@����!�u�.t��Q�߄��F9Pb�)��{�|��Ui����v�V��&��3ٙyk皿�,�T�+P��f��h��尯`�
߳�/9��Y��T�QQi:t��t�R����J�D�FP@z���4���.$R�I���K )�%|�������9���^k����$���ah>%~�`z�81�Zky�mCb�S�A"�&��Q�}��X�s�B���c:da6�;'���	仁r&_�mtZ i��y�R��tz�oyNocNCE �����N�����qˮ�.Q�2K��f���wXL�$�/���(	����fs�ly����nN���f��~��wVw�3V�_T��$Fj(㽰�F�}m�/era�؉�e�iٝy.�ͽ�]ߜ�nU��Tjr*�;�poS{�ݑ�,�w��o��L��>���������}󻚝�E=~���ۣ Z�Ƴ�?�[�	� {Չ����P�v��w�l�e?�Z�B��/dKҺ�����q�3%G>�6Ȓ��-z�7��˔����������tlv��M���I<m[R��=����o�k��K�O����'L�z9+dO��o8H�.�3ջ�z��=9�� �읭�C)���d�5l�Md��UC��h`I���?�}��Pt���z��R�#�:'�1HU�[�����"�zI�xZ��K0�	�:�zݔ$]N���A�?��kj���=�K3DP�9kgae�'�<��#�t�}��6�@^�\ǵة\4�?Z����M�G40��mLU�koP�W�X�2���.m��ՅJ�o���U��	� �1"y��׋���?�j}�!�K�\^���BZ�4���� ��Y�>F�m<���u]��<ژ_G�����;x٫//
�uxt�4�M�7}����0�Y!@�yc�Vrd�~i������_��kpEs(̭r~~K��Y�sW_�����{���f^xBK�(�e�[r-��� VP�fbt��ѩO�]���
'
K���Ej�k��#}�>$f� ��F E\��lz���6��|�Ҋ���������l/U�\�NC{{��a�5ϛ<����n|%������$���"_�|UsW@���[�z��>��X©P���`��M��ȫ� :�#��'��o^�	�Ni���at]քpw �/!�L�z4}��oQ�O�C��e�5Wia����A��n�Pś7 �� 󰽠gD��b{�A+X�k̎�*���N
��C��=!��˦�b~�$������5���߆���9Z���ё m�ٌ�[X
�������gՏ�`��<�M	�:DA�-�N�7q.�� Ct�\[�����!�z��m*v�T<|N{��7=֓�ڔ�Jo*����!x����E��[��~F�d�t=RV(;�!���:���D7���j�<*	���Y؞A{d�8�R�~�pu����hQg$�iP�椞
		�X�G��
��L�b0y��-��fZ�]�c��7�e�e���ʓ���̲ԯ�K�z�)��R�%oٖٴ��#?�U,���o>���.�Q�W�K��������@Q�5�X-�\�ǲƵ40�]�R�s��,��4A��IC�� ���~G�������4Z�}���PM�:#p8�R���gb���F��?��oԤ-
���M�O���Z�X4��I�g:+��ku���V��(��[�M���Wy&��y��I��_��~��:&����R��n��u������j������Y�/�m��>=�6;��������+}�����i�u�^W�A�����4��Ѣ3玮(pe?Z'�u�-Ę�E�o�&&��BzA\Q./7�>�Q��%����΢���i@f{������7N4#Z�Sϐ�;��;���O�����DJ�?D�-X;���u��3�U���E=^N��P�j��'�g(ex��s��P�����@���L�/v>J���[D.�� <�X��I��b��̔%uH�S4A��-�@�;{���L�8��}'���I�����a&��()��+��.#N�࣏!�4�a�/H��d��j�L�+�JIg�*4t�0_dg���
��˂��9 �
5Mf�+E����=J}g�	��0��)�X��o��7�9Eu�eF5>t�������w��f�c�Iz�.躙�)��r����P�C���^0�����a~���x��pÉ���A���<A�[��'}`x����V�:y��n0/��5O�(�(Y���2�I`\�)���Oc�O���-�����⫱��,�!�~-v�h����3���h�_�|7 ���������7�`����}��л,��P��et>�IyK�11	3�rd��$�h3Lr�`�R���у�i��/�M	|{3�˳�������{S��9bO�Ob3���������&,o���Q;�Xqgv��A-/��~.�����F+5��l�k⽬����9/����Q
8�D������K�w����ţY�ާ~h�ʲ�(]�t�#�j�M3�Gދ΅sz���nM4�C�(\��;R��U�C��J�µ�tI�@1���hv�id��@��/�����ε�?_����Ӝ�n��#:5�g�^j��`V����eJw�� q��9,�M�r��}�yg�Tz�D3����w���N���e���۝����O���xa��Pe���<O���zD=[�e�S8t�`a��W(���j�q�z�4��B�f�L�&��J�֨�M"O���������J���A��[�o���K d@[���>T>|�f�%Y]?Kp�ZX+�-3 i�d`�\/i�\��*I�,�B��lG��	�{5�6k�WM����Q�'�(N�omW�X���_��Ԃ��5(Ri5�#��'V�?Ӵ\t�L.F�`Lۋ'zObRG��m�� �O��b�aԷ�������E�������s2!�"��Q4d�i�;"�^n�Ô�[i ��5=��p������dyI>kH,hKC�rڨR?�[����A��_�$J����L�&��P�Z2�Q,-������x�?TRx"��<�PTFwƽ�����?���,ZoC۲j��<�4���Eut�C�Z��?)IU�/�y�]����������8��[hlbR�%�j^v�� �W�c�:�^wnѥK�1|�N�{����THNb/>�E���n���p��i��W���؉��)�K�'W�[��v�GB8Ll����|��$]�2UP�����1Ǐ3*�3�wF\e7VZY�i�\���I� /�؉��@6���Qh����b���b��/C�ge���Uװmt����<��_P��+��b�{����0w/���oBL�w����
���f�U]��f輯�����BY�t��t��9[�� f�i���q�A,��w�УB~Ě��S��ƚ���޻ /��C�l�8輸� =� ��Ј�!D\J��*���TskQѤ�#
��X��t��Q܉����F,k3�T�W�0�D*��;� ��R���Q^���lʌ�@���_�!D	ǰ]��(ƲFF�B�u���;@�e�����*�s"�)c�'j�'R�2�f"v����Q=�Xg������'�����i16(�:���`��2
ڷf��Y���m��D	�ӎqNk����~:���r�����̪� ��>Ua/����d<�Rc���H4Bv��0�	�:�����؇��h�w�6=�>ZP�o���ਫ���,��sD����wg�S�`�U���_�W���$/��nx_^]g�s>��M]��@���bI\gQ'��,X�An��!)e	���x�.)���IN�ҙ�����5_�h:�
��5�g�M��J-���\u�t��*O���T�M�&~�K5�$r��} �T�A����@�j���Z����}��zNt�>����e�z#	���Z9e9�Y�]���N}��ÓL����u�	P��8���q>�?����nq����N��m�/��m��KK��0��C������1:�0�*`�8�JI��c��d�R���GZ�J�� �/������}����[�GY'@��������]�?�q?Ò^��T	�e���;��B6�\���2c�a��$�osA���x �Vs��`�3d#����)J��
5Q��_�S�bKt��s-���Y�,c-���'	?�Y)�z*���;~O��U��.�=�>��-�0�o�U_6e+(o����������j���J 1�[;�C�6J��I��;�b/U��M��fn�y�)h�8�)��GsU�b(�I�z���wO0���#��>��0��:�1�d
�QVo���<��J��0�?td���J1g�J��3~�^�Pzp[r,a��o�H��0��|�xM��Q���'+�d�Dae��w��Éw֙��S\��3�Bb���t���=	� �e�R:����[��0X��,����&��:�4��_>�ϴ1��+~���������-{���\�^}��%������a�;[q�Mާ��f��**�a�?EQ:V��@�gvg 	�'" ��~(#���yE/9?�t�t4��sW��I��(OP��,�Șڵ��9�c����h���X&Jd��7hꮻ���;�w���7-�{7�NU5��?�h�;ƃ�C�ט)�"�?\��.��o���+9"��x3�-p�e�P[+2w����Xǥ�EE�I�þ�Y��ׅ~j��3|m^C%/�������r}b{��鍛-�X�������@B�}��)U��j����
��~r�9;=s�L�Q
��}�P��p4�&��/6>y��
p����vX�"YD�Z�=�'P���WecT�.c�6g�zyE���\?ۺ�-jKVL��܋��W��:�w�H�?�w�u^"�xj�9e����+92O{t���sAa���+����gT�G)��~ "�t(��|~l�,���-D����W�v��M�Ã� ͋�u�e�k����	Ը�Gt���#m����[ya��6��K�!
AΜ�yNl5��R��E+-k���q�	��0��",F�o������3	$w���ZX?ؑ\�L.�v䎒��Q�;N��ʕ]�1[5kx.���~45�Z�-@8�r�/��o�u�A�����)\�e�٩.�d?�$��jO�!��v�;5
v�3��|�!����h�.KP@e�ak��Y0�3��y��dd/��=�|~�h"y����*�Y���5���ws���QY]TX��zC��m�[��V�tUO�8����fR�Dʹo9���O�	FH����`����[3�S�e�V���LQR�L �{����2i皩�cv�6C�'����{K�ۻ�u����U��l� ��U���,��{��XcO�~�!��!
!�D�H��խ�*P�Y{0�T+��K�zGO~����J�����n����K��&��o�bE@@/�
�a(�Ms JDw���%��z��M#��a�g��٫1C��+s�"{Zjy������O����
{C��${>�0�n��+]Yx��D���0�� C�Nkɦwd�Sr����:(DU�*����.O^���u�$ئ��Hs�A���&�b�_q��\��x9Y������?7����F��k�NlK�$`H�BRv��i���Iِ�t�~L|��o���Xߚ-�bj����r̱x.Q�R⚬�辡Ŧ)QH%�cY-�W�n��c%A��]�)d��p��_��9��#�{���1�uB��j^9�+?��g�wiP�M��	f�C]!9�'>�9+����[��S4I���VJ��˖̳T
옓�E��0[��G�Zԉ%N��yib�gG]�ǈ�-�Z��E'tT}�(�P��p�s^;���R�&*{���ÖV�y�����V�Iנr�FF��8��-d�:n��K�� ��^����>��ত-��9���7&16>y� ¯��P�5]x���ٵ �}�k����vRH��͜}�9P�/G��	�l�:<T=Φ���ߜ�h�������R�Q���3PR�E��kU�#��/��:���@6�c=�RO�q76�K�$_�U�"�U���L:(�6,�'	��s�[K)���JOJ�a4('K�E�b��2������
�£� ���lcR߉w�HH:�T�^�4�)�|}T{\��>\�ys�l��5�qF�SpW�%�f�['Q'3����$ϲ����'ӷQkQ\�6< xْɁRw*�A8���\;p�zy�D 053)�e��2����h
Y����B�G�?���Pa)��zP�Č�_t��N��ݚ�PlJ��*��p^�P���c�'� .����Ue�3�Q�k��2�I��V�5ڥ^v6w�z�r��;��v©������Gɑ>_��������M�)�j�o�����ܚ+���O)|��}����5I��(�xb)�@B ��L�p��,��r��.V^��0���+�am�݉x*������{n�F�߲��)E�\B���Ⱥ�>=��+ɛ�I�t F!���,�����8^a����̖�iϠ+\Ps�I�l���%6zA�45�N��2��#������-5J@SuH'�Y��B�vy�Z�+!
��@���oe�[�e���)�����h[�D�Џ��,���)�'�	{�'4g��]�1�i�ΙSAE��	~�x����DV����U���`�PjU�y���P?�� <��5о�9��?�؝��95��Ѳ#K9��-�&�����\�y�β�=~>��~��4�7�(-ǩ�q�9�f��[��^�e=����b�,<�����1Q�U�3�����̓i��(52��/f�_k��?cf&��y�Ƨu@��I��l0��oJ �������i�Xf�E֡+��V^�ᤗ+*���)m�@Ŗqmƪ����v�7ր$�B�S�}\l�RА
�ͽ�~8h��w�v�bo�m�w��n=���
�{���?�7�j��qG&Z��s-�S_�1���ǽ_��Dz�E�EA�V7+<H[��9v�l��
�f ըV��i�s:_�e���N�<��w�X�ǽ��j���A�֜.t���OposS*ң�y~��;���e��sV�6�țՆ�=�O�	�fB��l�d�����{K��C����� ���gƺ3���2]cV��Y�N8�D���>���W�n����)[��2�.A]��#)v�����
��/��=0lE�3})Hi�GDPLh/@�|�x�.���I��IFgA�X�����`�SE�=�U�Fy�qؙF�u;��}��}�L����P��PV�H�)�}=J���_���*��4Kɋ�B��^�+{Y^R/��[E��Z��Fl������d�,�'�w����2���ki��,P��w��6*$��#�i$*q)"���z�?[X���&�S2�%~�{غ��KI61�n�6wV��������.�����V[7ބ�f��E�	@�қ��!��Lg�?!uPG���di�q��o�AS@;3�Hac/g:$z��r�ϻ�����$~X������(�n���V�gp�H�(��3�
j��
��AG��ӄ}�XpEG�L�E���=��&��T<�iX�!��	EA����.d-l�^e�z6H�.
�[���o��U��2�/���@���F�n�>����4��K��8f�2�s�=�VY����i�KA�C ��ӥ��7��Q3aSR�c���
0&O4V�q�� D߄ڜ�����*��������ד ���Е�:5�����2��j�BP��KΣ����;[oR���'�uzԦ�͚��(u2fG���q	�EX<��{Z��� �j�e�G�.% ��Iv����;ң"XH����h[�e֝1�tk�S�p�::�ߪ?�X[�)od��_߅&Ph����6�m�#�[!����Xhp]n��^�%V���Gx�ᶽ�_-���.p%6�ڢ����p���i�S�V���[:�	\s駷X=�)�J?jQ�5�� ��\��1��
��#\�b��qɠ��Y���d0-���X�߂~�5a����̭��M��1���NvQ��ٿ~�9 �ײ�;,�%�i-��
j�u�bs2��ٶ�v�O���d��O(���?��kl{3U5�p5�]0����T��|Cgr�=��{�JƦ��{:r��˪��ݹ�i�)h�}́x��EY��0���zǎ�L��%Yc���_[]��p��%<��0%:�+��V]��/}�!�G5Z��i��N�x�`�9�#w��Y�d�	�'6���7p,����;���jɴ�T�v�y5	��̪�	�qăE���h �����]��� i����=_Y��"��T>�%?�v�Wm3��c�fb 񯓎�����������0�d`m�f��k�������H$'��Gc�g�u��Y��iOj��ɻ�#}Z4�%�>o��M�R��71õ#�A����-@d����	���-���&��t:'����2�[�I?��grd��o=��H���Z��ђ���h��K����E�0�7�$+�4��E�-V ���~:.W�2x���	u�������u�%4�
���)M�ΥQ�'lv�)s��ƻ%d�l�hsL��=&:m=��������}�&�->bxL�bטC�jNH�kvώ���+�_+)����c�QZ�=N� 9�!�8M������������v�#\�%+o�����8k�ԩIq�R��A��A<1�=�9�b�*k&����G^�N����������fV:��{L����@F������'z��­p`J���9_�N�]w}m��|��7[~Wa��W5��2&��GU��|�/{q�Y3_* �g�`��'��>Q��nVv[���t(O�%:�i:1�S�߮��N�	�����8�
��X򧝯1$��\�5��lk�����}���_���q@�ݦ���A�oQ����� �2=��S`v0]��;�3L0��6�x �A�R�Y`�d��3>�A�|��7��3��%��1h��:��kwxBk�ѿ��Z��+x�3������lp�Nd���24#�x�]�Ɇ�6Y��D�T�pl�E�{��d�Z'b���������;z��T\��ʻ�'��?� 0a^�eA���Uh�O��4�3����`k��{�9�Ԗ�q_jF�� �2'�
�%�'�Td��jE�|F駟wm8��7��~R���ʞ�㑺r���Ɔ-�����~���|���M�-M'Kk�M�0��ޘ���z�WN���HW�瓝�K}gn��<�k���~�.������u��O�����XoZ�'�^@cG�J4A��!���-��j��N��A?oɣ�ki(�32��9_�y��O"M$�*	����񯙓&�Y}���qKͫ��2����pz��+%,7�����$hv�׹���e�A�%�;�*���!D�z�y�
LX������k���l>/.7苅���=MQ5���E�U���_����+��^tԜ�L�G��K��uy:7�?(ނuE�D)��5f�v�ǉ}��J���t���5�ܑp���[�vhe���M5wr�Xo�O�����'�9���'J��d���Z�j���ߑ_��s����̍wP�)p�V��.E`����'o�'d�����Չ��O��+M�_��v�	z�Aw!�g�ȋC&4�v�Ž���U�tq�sЗa�� MM������ms��<5M�c^O��=�ePg�ԝM�֟�3�T%���ى>�gA;r����_��oX��}Ŧ$��γK��xC	;B�h��9(�������}�/a,	g�)��(�(BW=w��ظA�D'9�ĜOwN�۪?Z���tG���L�h���갲��C7��[���Z���+*�%ɳ��+{U?�UW5�M5Oa�/�`//*�X�+z#��!8K�έ�1�j.{%.ٖ�x��܃l��F��z���#H��Q�~�56��.L����jD����l�Bu[�<�~��
���!D�T��\�g�tl͏�>^^2��2��Cᅁ�Y�r��@�Upߵ5�ݏM�l���(���c|ݧP}�
ԶG�@�X��M���W�waH�Eɷ��Ϊ�x��"]�N�~�i��	J�|�@.��N�"�=�mM0�nk^�����^�^<\ �a��O�_�Y"�����?� @q��ٽ��Y��**�9��b&��z*��nL�t`�@�{8�沝�?/����?��8�I�J<�1�A�\��
�J��6�k5�`*�t#��6���|n}}��I�5�����|�7����>��$��&(Qu�a��uh+h��=I�Ϙޠ�!�|
�oR.�B-�Q�C:-�C5 �r��WJ��=�d�*(����u%�Έ[7�շ�r�7P�0G���f\j��q��+�����keI���=u$]t@�h��
�X��b�����ݘ�ɝ>��g2���k����|3H�ZrE��1��c��߆WK����h���H���c"䌧�q!�)η��t�'��P^l�Z���R.ն�>O�F:��??����AKy�M�6��B��^��?-��n�$*:��L ؐ�yd����vA��#��,��i�D��f)�{Sv �k^a{�T6��V!�VGp��b���]\Й,?'p���=l��w{[�.c�Z��1��^K��"�tt/tQYWʍΦ�I��M�p�/H���!&�m�lg�'�"	����+� �:���F\���c[n����n[>�Q�\:u�5c�
��M~�N_h����|�?�F���an�\���N��ә�@P2?R�m�tx
&ٿ<��Bk)4�IOs��r@����:Jr!���Sk����$����������v�h����l�r�n�I�u�S��V��).��L��^��y�y���먨�*�Ç��$��~?Q�6�L�o+��A��H&�5�t����k�`'�u\D:h�u�l �z�� %J4J�u�����-pI��j֮��Ti��[���p�2�4�~D~�&b���Q �^?�:|�4:^����pL��Vq�ej�� !���03���z�������A#]��^'�\�.J ����|0�ͤJ�p����'{|`�7�H^=�4&�?.�p=�P��m{��t�-u���$�/{�{��j	�O��6�+b&L�S��Z�92�,2��Y-�b ��p'�����}FX�9��'?��qF�(�c_)�`�:y�#�^�A�8^�;y��
T�F�UX�]�@ �n��cVҗP��)u��4��:B���0y7��H��~�l{��U'ׁ��!�p(�{��UNI�i�ڟ���T��y2M�#�(D^���/�z��柘9�&b���Cמ���jo�$&��mN����)�Z˃J��������Zd����]"�A�q���fW��:s1	lÒhe��	�[�i�ʖn� b��:��F���XxV�F�*��3��g]^��rX�l�MdQ�����voU��w\�����Bo]��sVU6t����� �)/R
㩨@�0�dd �Y��e�f"�4���{Y0�h(f����m�]��ԥ�Bm��B�V��$�G�#��&��9���2�0ݸ�Ǣ�f ��׹�W��ֿ���G�L�%�]��d��G���7�����T :*�b�q}�.tfV�R�%鑝;%q �vzKw�۰=r�W��@�d1�U�n�!�V8\�K��P�S�����y�z�#{\�0���8پ!��]�&r�ӓ�0�1����B��
s���E�#�\�LU�dʲ��vܱf�:-uHBA�O��Ti�5��`�G1����}R�.\2�Sn��j�Bz�U�m9��_���A�n��B�#���p���������*y���"2��8�AF�Ic����_=;}�{fe����*'k���$odU!,!96���~x�o�T�����J؏-���~1��q:��5lվW"5���I�������%˝�5֕&���]|)��%�c�-%ک��I�X�纶��$�:�f�t��($:�v-
�N�d3�^�9h݋3�W+\�ؽ9��<��s���7^3,�]�ai*S'#1�	�����;�.�h���c(&��c��� ���ّ�Ed�!q�o#9g^�}��>p4HI�0�C�l�gK]����������o�Ő8c��S�l�In�=�[�gh��k�(�iV ���?8��@�Κ��{vƏ�o�.�|�����	��	Ҫ:�����j�2��x�[Ԣl�����j1[���W�����X��k8��mޥ�^:��EhQ��/D45`.�$+���d�L{�a��|va���yU��`=��x��$����2�z� � �	�Y��%�#��6�ug�j�ͦ$���`�b���g�3f��\qQU��V7�Y{>�5�oHU�]� o��e�h�����5�h�z҇���s��_��9<�c��9� ��H��[Ma*%�Sccr�GH�^EԿ���=��s��>���M�w�� �Ap�j���'�����ޫ�ݸ4�,�	�N�T(����%���c��k��t ���M�U˷:���49˖�ǡd5��@��)�J;���?�J ݗ��'y��B��u��]��r���-���p fQ�UȦ���A+�Z�jXi�I;� 8�]Tn�Wt�J1�1���b��^�g�D�7��[,�S����!59��$���"��}ش�Ŷe0���\n"�H�|���XzS}�^���$ɝ''?�II������8��R��,S������(kÝ�
+|�Vk�Z��!Q��T���,R���V@>1�ΐ~��[.t�Zx/�/Á���������D`�w�3���n_�w��x�p".�Ua���׃�lY�Å�n��-�����x�x�d"w4~Z������iT�˃o�uS@gu�#1N�{�ȁ��Cꄳ�C,NP̘�Cαrs
�D��j���4��j%��χA/Ӏ�-�@��Y��UB#�[�XG��f�����.A�yA	��웱����by�Dv�Ļ�*_���LsSs�WA�(��'�><����kY�pS�Ę�
>/��Gi�֢=���-�Ŝp �ZK�.#���LS��J�+Ie��g����� �a���5oyS»q�� rd��<	z��k��ˋ�}WҶ2&~@�W T��re�qG���%m�=��\�-9sd���.P� Օ����ݖ��˩���m��(`�A�7#���(���Ts�+����Ӡ����i'��%��_��\c�	�u��z?|pMb �{��|dgQ1��n�S�U�6�y�͡�KY���v�N>G"���W�^�0;!��[K^�]KlT*�$Q�z�O�Fl�5<)\1P�s(.�w���[8�Z���t�e���R���Ԯ�`w'#�,q����g��t��V?�4-�f��kr��NOP	��Vk�NP���(S"��pP�t%)L��Ȋ�&��d�'��}��7g+�Z�r���6��.B<t�ZS�\8k�9C�#�`G;���e��S��*�̇ug�d���TS�h�BL�Y0�'�3����KE�P7=XJe/��O��)���c���`����J��83�j�>��[9�M���]}�����﷒Fu�n�oap�Qԗ5A;��ih�Bm��{K��sU��<_�������X��V1
���Oj�7h�����plݛ:����Gm�n3'�ř�;�������k�j���y�g�`~d�*e����2UU��X�ޥ���(6��Nl�Ru�����c�鰙����,3�ga#��+�;��y�z���,0#�;O���ظe�L�Pp��[�v천ZX��lZ1`�@����;�!z��6\�6/J�c�@}+D隷�S3\�ރ�*��m�5��:J7�a��f�*��Y��۱�O\�:��绂�F��v��Ƶ�з��=`�#��|j��}i�l�ٰ��������r�����o �%|�� aw���f�&��ޠ�6�hԧ³<Et3{�䩅cej]tw�}��ݗ6�߁�O���	l����G�H��) �yx�:ha6�q���p�/Џx�ti����%�+C�㯝�RҰL��<��ԑݣ����3Ml:���*���ö(^��.(������_A���)x�����j��F��;����s��?���zg��R�0��d/δ�K��ޏ�� ��$�`i���=@}4��wBӔ��;�3]��uڥ�{a��>���(��`źϘ~��44��`�l L��-�$ @4�G^m0�	�?{pf�eZo��W0��:Tc�)3��RI�V�t���ã���.�:O��$P(��l��p%&{P	�$�X�h��O�h�����:,}=��\($Sf����4���ͱg�Mu���Y�Z�
�B\_���a�R�T�����C�>[���;S�.Â{M�����@ն�D`�#@!6&���^�ٟq��E��L|g��u�������G�m�#w긁����t~7>*��"�!�C�J�٠5�h�e"�d���u��nZ�P[���(Q��7�e�R"Oq9y��h)=.3��X�j���VaVCO,a��@�U��1����FW�~�fml����, y���\"����*/s�`@��?�����~���Ğ��E�l��5��i��y_�Z�[�[�Q{��i�`p�%�,��k��O�'�b�?�����m*�3���4�P��px�-cB�`�C%Y7��P.�6d���ii�d��Xa�j"f{.�2*�\�l!zl�@p�шPdȐ~��2U����d����+�r+\��J�7�'R�ɬ7# �ԅ���B� 3x�arwTF?�_u���3�5,��]���0��(_�V���l5&d�G>l"�#��~T�q���x���^5�x�n���m���Ym����rhu�r��h+�6�.��u���~ؿG%`=l���ƃ$VpE`X�r�6ݠ*N1K�h|�YV"[�U1���� ~5�~��G�T���;�;�o��Ȑi!$�Br�n��ka"�x,�u
��o�V����㋼A�!�bh�9�K���,����F-Dsv���@�?�a9�`a�[n�A�A+��������[�.K���$y`���T�RFD�8�a��:��瓅���'�ٰik\�y�ߴ���B���N�]�ĺӃ_�T��	��np���*^~�]�^hL���z�K��P�5��E_��8�!J#]�#%��Ŀ�Y
Ԕ�&A'�z~%��$���9�I5���zHt��Ϙ�b���)��%�G
]x���/|���Dfe�m�c��0x�jbx��<!��D�p�+z8h�$2��Cbh��@H� ɟ�޷�íd3"Τ�'��*z�:v�e��:����]��^�z��Bvu���(C��pF�*��d��*(s4��?;�	̅����Td����iNM��K��9��жTn	L��mY��
�L����)n�2��]y�T�׮S��(�h���#�m���[t0Iş�\��3XG<S���rRxI�^���.A��v�Md��]f�|�z%�3F��k(z�����q�D�-�nS�_e�]���D#�����-��o�{;����7,0����E���# ����!J�Wy�����
��'Bx�E�H>JC�d}�U݋��B\xۊ�SAPJ��FD�I�/�`r�5�.t�<��o��{�f���6	_빺H&�t�di,�L�V,���$�R���J�#r�P��Ece�6����LdW(:Ȁ<sj�:H�-�E�����������G��}'ipJ�WĻAS�k3Љ;��>�/���i9�;����~�_�e�7��T����e���Ag�Zz��C;�����U���Ȕ��|u�me|�r,���ɼ+��b�R���>��@PP䫣TM�X�>%� )p�&��[$�����bH��|���L� ���0��@940���t�e#���0���W�޴;�b�)n@C-�F�Zg�i����I��W� �ݘ�~�&��)1Zn0[D��L`��|�H��נD�� ��t�!W�l����*W%/ J+�~�������(�{j��z��}Q	p��ow �Z� '�33�`���FYafZb�[�)�5�ٺh��SB��"^�9%R��T��j�j'R:��l�D�c��(Q���������!4:�g����Z�� �2�\����:9�&��MGJ�&�j#��T��w%>�KW0�.��6|�h���?�O�P�&���֭]��~
���m���jP2Y�g �y�mn.��d=�`�]}
�S���5�_�#�ZX��΂U�֟cM�K���3u�'��{���֌fb��SnZ���[�=V ����d=,M���Æ1��pGȐ�)�x�e�4�њ��{�W�w�\�ϳ%��5���w7E���,2r*ѪE�m��l�d��rc�Ѱ��?��:n�I�z�����Lf��Y�ގ(�\�W�9��gU
��J&<�׮F�S�#Ug0�6�\3��YN�/�~u �"�d�`��SC�s�;����.�̺Ш��U��xS�h�\�H|^��^��޲�q��EYU�G����iN0Z�9��d����;
n���!��-�����Y;���ZN�b�˞������~F��+kpWB�m�o�`�� Q&m}�x����6�ݖ�h�^O�������}%�(�@�j��V�"t#ҟ(��f���0�(�r�dQ3�'��@䕧��U������|�y �-DΣ�te�E"'��K�%�/�af����z�ϛ~#$�!T9_�`�P8�i��r����)�XZ�8�8~H}�DR+l�yj�t=��˘�t�eg(]P����B��-��\��G���+̪���y��yǯգ�-lG	��Ô��U 	�B'��a��Ma1���'��'+LM~�3a�Kqw����%�3�����Ǒ
��ҧh`6'�`6��:?`
�Q%�������xXn
�� �����C
�&���n���JR̈́>dc��7��-eo-͏�n���5[���c�s�2��E�'C��ȏ��{2��EF�
�O٢��ږ���h�y��w�c�_��v���̢�5))��U�ɺ�6$����XM|�m_�L�/9�%�>�ɼeN�cr���w	o*úL�!d?��>�қ�z8���� t����W�@cQ�z��\_i�q�wj�.�[���t��8�>�BpdXsX���B�OV������sv�D>j��M)2*%#�:�Jb<��%@���ٲ�v��Ւ�v�у���/7���98����ߺ)XL�^;����� s�:ȧ���	�/!6-V�@�\v�z�ޕ��͂k��o˨� ��jD*b���vߙ6����P$�w�Q�A��ڻ��:KE,����hn�)YF+Y�]����ɴLG�6�N�չ���qth]Om�E�=������R��s9��1?b�)f�T�c��vy|�W3v�a7g���K�W��$�[�>ls��@�FCLE�#dlP�&_��27Z c��YH��8O������W���W;����f�v=���X��D����b|����u;Ѻi~�Z��R�n�ќ��V*,��g�꠲7)�3t6�����	��k�o�_-��~tR�h<�v�A�����'�	>�ڵ�}�g¥��~�~��X�<���ڙ�\�?.�r@a)Spٺ��#���\��񑢓��"B�NI����rt({ٳGQ����RYRɒE�=�n��,��>�샱o��{F������龯�u�^����|]�}߳��E�jVb@���'��=��q;���$=# ���̉�vLk��evy�h*`0�O8�g����6I�S�|���q�ļVK�6I�0���i��^a�ޭ����?NRʱ���	�����
��4.�0�7�&�k�:ה�T���z��қPC��tJ������x>��>�-���G��l�?����M#���.��"V����v+�۳���� O�+�x������1��ex��j��4a�Fe�������)G!�Ѷf	���:�v����!G�w̶p.S�K?M� �Q���"��@�_/��`�c"�\���ETje5�fs����?���KA�L��P�Dټ���/��q�t�餧�}~���E���~ �
Ц�� D��f�o�MI�/z<W�������Z�I��̲f�y�eT���lwΖ'eF��!�>�T���6w�N7����_�u����^�q+'�|�����`"\��:�9�������0KO����n�E���y7��u��v��S?iju�z��KL�^�y�z�v�Qc����l|cOu)��0�'��92:|����ޗ��S.QW�ٌ��L�.JT�Ga�/�[�A៩~�v�ZP�1宫>�[�3�,�H����ּǵ��1t���`Ƴ���
i��� ��c�Hy��{�� &�O46j@#�{!���9=̧<
�2}��9�>Lw�=j�R�Ҥ ��a�2�M]�G5�\>g&n�`��(p��.PO�o{9宽�c�Շ'A|��/���/#��E�f�$���β�?}.��n���l��)��GYK�-�G�dzKΣX���#R^��?4��j^a���u�b�ř���J�v�O>-���_�̒���j�L��S6��+r�:X"�!�5旑���Gj��wG.�t3\�����{5R���ܞK_�-B�&;Vg+�a�3U���hk�r�e�2�Y29aP���z�3���N�*�4��Ԟr� Z�$�q��c������%�6�s[��ɭ.�s�4�o�o�;�~�ϳuD.��Q(`K���+����.�%�Tunvx�T�'4�A�d�c��<��H���S�-{���j���e��<������^�}t?#c��n(�?m�G�QG��^��Cv~r;��Y�����N�E���I)�3��r�<υzS����A�_ab~����W�5h�t)�7�����~��2;�����%rȖiF")#֡��'�+[��Ҡm��j�ԙ6F����\z�_�F޲��-*��!EUBB�\��,e�^�wi7�ps1�O}���B�+4�?�a���Cآ�Y�X�_�2w �Q�3�Щqk�B����Ϛ���\y��&e�=�C>�m!���+�a櫕�zC����6�c��9>��`��u,ci0��ު�Sm�c���O�JwNk�	?``�7^Έ�\�;:��H*�k��ut�H!7�F7�ӕ��7�QS��V`�R��^�:��,���cH�g;��_�L޲M���;����`�y�f�߯m |��j�8� ���������c��Ģ�a�)<�'�N������ ��w�Gn�D���O?��U�Ö36��DM��B;b�,����=�m��td6�R-Â�3]ꮏ]Γ�y�W0��I�P�V�'��S�A �O(t�5�m�+w_��*�,��[1%�M��Ѝ�_Ɍ�@�8��c�(XϕGH�A�����8���@qN�w�c�i���%D�PU����
HJE_n%o�-����+��w�@�) [@GD�%�N��u.��R���.��µ��E��s1���Y�K��MN��`���3[N�W�(�S���w�H^wד݊��]j?��J�ln��K��(�Q�jU��m�ݕ�1���h���������X�09�ݗ�d�C(�=���[&%3lw0��l�"�����ur���7l����߹�c��|���(>��S�T�#ڮ�n�n[���n1�CrG�*f�j�8�.8���5���b}�8o�/���%��_݈R�6�L&��2ϼ'�R�2,�Xr��f�l�cҎ�S�%J5w/��Y�2;�[e�q���5-~H[T�㿟@�csP'�|����:|�͝�]x�A�k��CfԂ�3�W+Z�
��/��ܓp�M����om�=C)��(t�AD��O�<�U)#���lE6�p���/0��(X,��Ŗ���7��kn�q�z�� �`;E�+���;�������*�5mvc�
�!��&D�cu�r�/�SID��ݼ�Q�߷�׹>��U��F��'��?���$�z����[_����m��s~#�5ɋ�e3,�%��5��q�A���k5`p�� C/uq-S�oѨ�_G�e̯_�7�F�Z�/E�Ǣ:�~B`E�}R�I0�5�E��?�ڑ��Zj�wɻn�Av	��a��g���y��Su�f�^Bgz[@�Q�����2:I���i�k,�|0	/����1�8�����4��M�}�r�Y+�U�C����(�� �^5�������7�P��x6f|@�n�L��j�F��龃q�����+�-=J$�ti�:��Gh��k�$>'i�D��.�n�����ޖ���R(=��˭:��Y��6���Ȗb�!8ws�����#��`����Ʌ��͗7l*�gq^i���X]�b;�ǵ���2 N����+�3b��J:/�Y�8�`��0ܥj��hG}�(�ϋ��r��4�
D�� @Y�	�zˑM�ۉg�`����܄��ϴ��Νp�\e)

A(���Rs��xy�w�V}��x�6+de��LA�E]��b�V�<�׏��X$��fͫ�u�t=k�jϽa���7 �mnb���ڒ���wz�S$x���>giH���A�.�V\"t~C�\���e����'��%�2]q������SW*:��S6��U�5���-|H��or��_�.H�����
��E5Ϭ�����F��n.·^'d����zK��*��3��u�<�soAM˿=�g�: (�7��ߗ�/¹�X�-w�
#,A|#OEM����|�x�+�V�d��T�%���F����?Mi�Y��;�_��G�T����QVS+ܝRX$l�&���
�A��ԴV36�*x��G�_���_���TP7hud7����z橥��Xt�����Ոpa��-t�J4'k�26fo���V
��Tq�P| ��ss!|���`�+@��o:P��1W��9�� u�Ÿ��M+���-�}D��V"+@�	ـ��9`���o]2����߂�o��~6��K�X#�֬xJ��Aua�_�p��A<�Q(�@6���B�(��^�����Ÿ�e>c�>w0���?����K�Z��ѻ�v�K���<0��I%o�Yʮ:�$�vS?�L͍��0����ާ�7���$���t���t���S��Dg��գa��T�z��=]��K�����<,�ɬ<��ۏk'}�1�\n�J3���9�B��f������?<���Y�&h���H�Ǜ�b���Kݑ��֭�"�����١�.�����ذ��p�qWש���w̫�ӿ��7�����}t�RJ9�E�C�M�C�>^@����-`�)og9�`����W���g�@�n�pd�ޕXɱu��=�;��3�/s�ҹ4��Kqgh�����q0.��C�DK��~|K����G�7�_��8e1�Ov1���D�ׇ#�h�m��Z�5��GNF-dAo%�7��e��Dd�?�L�6����j0��ODy.��Z���
'�ۨ��1� Y��x�^P@�f��a�c�5n�H�_�$�m� ��,�Z���K=��Y�d�zc(I�k0N�������C��
c����B˩��W�˭�'�#����(�mV���T@��#���o�p;SQnc1���*v���W]�]���/s�����\Y�l�����������F��ㇳ� A���<M~�N�^�a�D�g�1S)t��e	�zJc�'��
W)[6ײ+=E�F�'D��vE+	������=M��������j���UR��;W�=�)�2�k4*�e�4ʂ��^D�VEF�f�?���1��9=\���h�ظ2j�Y]���J�\A��2.%��LL�\s(Y���}*ea���L-��=�_	�|�U�y�`x?Hu�./q��+���Z'+�I6Jo���!XB����i�Ն�����k�>M X�٣��4C��s� *>@��PWX��v3��Q2B*i����CD�bQ�� �p��RAi��(?2�x���K��U��#��4�m��ʁ�t��2����>	C^,�hh�b;'s�(@���������D9٠�N��.��z��=U���qVWB����h��҃b>����e����s�K/����洗��o=�v:��$v��wr&z�SJi6��\=��}�'�C��q������)|�����,���ۏGI�˻�}
���&��G�I#��,�����Dߖ��E#�o�#�#]1��y�2V��i�J�13xS.�A��g�Ұ��M��,�:���Ʉ�M�	���ȃ4�|؇AR�,O?�u�hkQ{� q�L����-�q�,׽�=/�jH �72��s1ȇ��dbV����f��T���ҹ�ֺW�@�e�4�;{޸t:�]s}634��p�ȫ����})��3 �"A�ܟ+_,�ה�>y�B�b���{��u��bj����~���&�(P�_����?�ʻL��8��kO���xZ���z����X����4�	>���​�&�1��NV�g�����2ͬv]��0r �&�%f���}`AR�,�r֧��>6��=,yW)U�fn�^$�*�zو��wB}|=�sAw�Y൏�8��Ct��8����ՠ�v�����\�w��﹗�>��l��#�_�����R%��1T�9���9y\���/���4�uKq�@����[�k�����Fs��}���|��JA��bV*5ũ(�5��;-��!;a��i�-~?���'B�1�\!o�s�69<�w���4�Z~׷��pާ�X�+�kx._wA�"Xk��I����5)~g@N<�+��kh=��1��)�e_j�2�y��K��A-����s�`�ݹ����	� @{� �� �{��$&��� ���5��:QLn5�G>�1Wo�yc�?E�c���p�hF��*\�����K�0r����R�y��v���R*���gy`����ē:��9�oB�#}�M&�щ;W&Ke��vJ0�.��6���P�7`�o�V���ɬ���R���2���~A{���T��"�>�J$&�ށl�g��@4)$&j��_"��h�!�A�kC}l��M@V����*�c*�U����*ZL�~*v��ZII8�`(k�����ޡ͑��AsP]������h���p���պQ.���-�Wqi�,�q]CWҒ OQ�^"_"�Dx�kw��,u�zD=���`����qX&�9����8�y���a�B��qB�:���U|��t���E��70@�e�(�9�S�a� �fG2U�l#��7>�9�����sEf�R˦�,�z�`��}� ��#�|��Ј�b��� �>eu9*��]Pv�wr��s����za��Z�z��P�WcYŌ���8�<p0c��N+:�LN�+v���g��g���Tmi�0^d�{3�Y��a�SL���I+�	�6,�]#��fI�'�o��d\��b8@/'GTV�&�6�'��0?!R8���Sf6��ٶ
�y�����[_��L���I=��Ȧ�B�'���(:Z�E~} �t�Y O�h֦z"C���̩_�����C/���X�+��!TCq�\640��z	�Qm���	+w�2\�޾}Sv�}4+�'�9O&R+7�W��7!P�+�r�'E��m�]%�ͻ 	I�k�v�\
.��B�F���	��E����aH���_\
�;�z��@,�������<n60]��~���p3'�/M2B&�_�=Ȟۨ-c��i40����w���=�FI�:���R)�\��{ݧn&�d�`�T�2|�}�O�>�*��߱�c-�O_������M� �:Y�����ά�8���tI�/���H�*��ĿM*eڞ�^E�_����cjFo��B����*��߾/Q�DJ� (�˺�l���^)�Lt�v�~�>��:E\��ƀ6z���x���b���`��T:��n	��U��2��A/�k!�5p�	\���m|������5jI�����B֕�]�ݟ5��$С@т��H�P���.e� H?d#��>�m{��}�K���ry��8�D�嫍OT�aG�$ř�+	��/�rB����gxh�6X�|�j���db�ξ��II��C�&Þh�� V�4-�j7V���7�����ů CB[;�F�%�Ȃ0ˊN�<���}�Ӵ�e}U�ؗ�6A�60[���}'�&��2��nN'A����#�e'�e����F���=�m��h���n���{�F�Zo����h�=��!�"�,��=�[��֤^޴)h�����E�1���3�k�*��[�m9T���}�g��ۀ޶h�w��7P���:/[���2���ֵ��X!��(��*��!�	BP���2޴~M�vxM�p#�8��W��^ؖ�����[����S�"т�qz$���j��O�?�-��3��̣�m�L�t��
],Xr�D�#*S�Tt ��!Y��lu�� f�~�²�Ke��+�>�,��"���Iqz�Ç��Y"�ȶԋ�=��j ���ҿ�������n�}�~Kp����߫l��M�+Y����d�kD�r�J�K�j�B.�HɯH9hD� ��7�����ؕ7�!QG����X3�h�Ek����so�/�8?�@�j�5�.�=�a�~.��2'ʹ�VIKM+�;�XX`��9Fj_�(�[�K�L7�(A�c���]��������q���Y�fr<��9" >���f[c9�������W��z(���)P^ +e���\����
0�F�ѵ�&~��0h8(?p�"Q���	ӸK>��2kv[�er�P]9P�E���bt�\n������8�L�9����˼G�4��� ��̓�^��w�Ӂ_���bS{���/�!T��Q@�({H_�m*0�}&�d�!\��2�o7�e�?����a3=�-q�$W�=��)�o+(�T�_n���htgV�I��4�p/�N��hdb���#��P�N�x�1�=������������Fs��bXz�����P_�n�K�_Sg�ꤵ��F�L�Y��t8�{�C�%��F���[��m���8uT'�̧D+=Z��'<ު*�Q�h����:�:x��f�oE�_7�3�F���m�����/��� �T��ܲ����Oc���<��%=0qU�64i�*�.��U��Z���OkRp��ı�c�֟ f��Oq���>L��J|ti��Hi%r@�BM%���q��#�S�e�\���(u�^ �n��>�{G�aVHd�ѻ��ب���Y���������4�=���Я-;������ʯ�M�A+Q��K���n�C���@��բ������J�Qf���I�9K���Ҳ�!.ݬ��ii���� ��.&̀��i�Q���2�%U\��_$m3�%.ޤ�H&��"(CnT�Y|"�}|�+��ÍGP'��S:���|l@�9��}��Oc�9�ٱH�:�g9U7�4�1\0j�.�����1��~����HL:]`��-��r�����h�C� dF��YK�n� �^#&�S~2#�H�@��S
"K�D�x7�FP���9o���혪�7�6?����nqP����@�z�|j��u��Ά$�$ ��˖� 2)#,��ihi�߃=������D�C#t�v�-m���;}UV������d�	*7}�V���@Gu���L�Ф�-Q`�3�PC�.¾�Z_����kU�7P���v�/�?����dYA�:	8����qF���	��`��*l{w+����Ä�ˍX$/�{�3��4Z�K�H���d�>̲%��_y2�TFJ����ͻ�nD�L\�y�%���ѭ�8����0����A�_� I�b�y���Q�Y�-Mu(��U�K�.���@�p�����L���SH���y�s�zg��?v�P!��1���+�PbCJ���B���1ɧ�s4�0�a�)w�w����Aփ�f�g��R������0�ˍ4D6_�+�l��x0�`��cNM���j�Yخ�a9;]���ϩ8j
̈�ݒ�uvD�>���[ίY\K�B�V�Ae-�g�8�A~R�H#���wV	H#��ns*�`�����/P��z25��vU%hUth�ߢ��5��K���@��h�����L�dl���~�F�>n|=�lA���n�""���~� ��٤�?�m�)b��~�r-�krI'��-F��r�z�E2��%[������cfv�֖A�~�kc7v+��-E�[���ܩW�ڶʉH//�-�O]�S��t���3�K"副^�ʣ	8�'�ћ����Y�Gp|�$��-ktڏ1�"���'�8@��aP~�*��p.���
� j�g"߁R%yjŬ�e�D�Q|�j�� AH��~��pA���Ud�2�y�ƕ䢲S�ܠ�W�q��U��}7�v�}�(�R-
/��uu�֠�ӏ�T.��&���uR񮸧5jLG/��<gY[�N��l�[�����p����B�ߍ'����t�t����nF���G��J"*�7�ɲw
�,����s�������ҵ.���2S���p�8�aL=X��^ʚ�*T��v3�u�nrlZz�����}��֊�E �4�3��&�7�6�a�'��hD���� %F��݂WWM+�L��:8	b��a��1�p��t��jL�u�8@����<��D�-����,��\!nCU\g�ˊ���n�����6?;z)G~k3�|R2N�����n�e�lnn��.	 �	����������bIx�zN�J)�l����	�y^�l�Ey]C��(<�׷8��"S|(R��T�c&�{?�eS[n���ԕ_,�E���A�Pޑ����.����(���:4bQܫ&�іp��ƪ�M���St,��e$�3�=��N2�J��[��&� x28K���y+h�roZJeg�{�� ?��+�t�}'�|�]��$���?��8�1���'8�ÿ�S�ڲ�������{����M)��e�m����T�	��i�W�"`���5/�ˎ�rzMGbvD���&��M1�B`�^
P�$̊� {��]�jr�������s魤�qs��Y�j$#Jp�{��~�.F��5�Ȇ�g�q}}/u��Y�3\ՇT��1{e;W�.�<8
)����w�V�P�:�n������G{b@/�1�� K�\.���7�Z�n����ś��8y:���IC^H���b���l��	�A��q���Go��d���=����W%���̬��ɑ���:"*�KY��/���I��.��A�����e��
-�(X&~4A��x�/ ��������I��E�5�IA=ݬu�c糼f�9�F�: �һl�Xv&�3���:�#���>�Jٳ����0���3b,��jg��N���̮e}g�HN:>p��C��Ⴣ]�?��Su�@�f8������̂�' |�^.ڂ~�ci%�����E��/��4��T��ڹ_}�͆���E��"�3J�\�
��&�����~�ř�X'���ZI�	��n���+~Bu����e�VdN���*'�+2.�9��(��󛻭�3��>ތgǦ���Xw�g ����k�F��8�ʤ��S'G�?��7����^���~klؖv�nǢo�I��La���ay�����8,��Rp�þtv�'<כ�B��7H�����D��A��Y{t���KX�2�t�a@���좠�3��� ��ۄ���~���� 3�K22t�䩿�֑������P�5�+��WR��N�*�(Q�O]{'��r�9&턵��i�I  a�J̨���/�O���ͷ)�5=��y:	���GV���G�`����é�WÇ�B6����P�V��4Aۚ^�V���:t�
�f!NO��y9ā��\�>8�̈�Χ
Ħ��DnE�׵1hm��T_򗗯;/�T�`Ķͭ24D>�Q�����S��%�k��
!J���.� ��&W�?�a�{��Sǎ꽠m�5|,��)/�} ����!!\_�i�����&�k�LE�C��Q4S���p(�������u=cg�*���5�@�j�u2��%8_&	'��E���U���������+x�H_�奢\��6f���=����Ow��R�[�`��L�L���������ja����X�0�Gٛ��t�}�����D@�_��~1c����4��w�p��R1�H6�P|9��ŷ9�:����
���2�1�)�vī�ߪ����^'����ö,�������ٻ�r���[sL��o��	��p�\���u��m�iz�<�KՇt`Y^�am�́�NhR$5����R����c�O���T��9Z���5Ȯ^�CqhI�Uh��ǌ&h)s��u|�ڠW���!%�U?'?b�a T��S59?�]�Z"*W�d�'�Z��JG��t����� ]� �t��ny"	��!h��`m�츇��x��N��境4k�,Y�EٺI��ub,;���?	�_�z�Bv��[:^��2K#�}!��X=lބ�����DKP���ڛd/�u����N��1MX�W".D�;A�|��z�z�>OM4��<�Is���,:S�m��e���M��^��Z�������p�4��?��o�2:g�@��QV���!�A���a*�H�EwYLJ*%J�%؅<2�ux�=�0�V����B�k�v-?x�L[��GW��uc8�V��IK?q�U�������>B`��r�o.�����7ސ�tI�[_҄Ž_�,���L%ORi�ut?b!�%xt�� �6��٭P����b喕�X[4:E����k$Mde�F���H�r�-���1M�da7�>#���vL �ی��z�gt����u�f��yc+���!��\[��"�
	�>iQ����H�Zx��LAZR+i� �1�o��S�Z����Az7��h�L�y*�D�}��R2X�$��j�߱�Dx�CN�5���障:��L(H�=���;:�`<3�QOc�,��ju��~d#g=b��E��(1���=���n_ �2�����=&ъ/{��
�v��%�ؓh�r�;���%�7˵��N4Z�H"��o����NB
m�M��` �]GЕ���wV�*�.uwll^5�yih�.���0X��\��9�l�~R�S�^��Kx;�!~$�ˠ⪇~%��9���d\	zT6���s;w,��
��E���#Q�|�f�T%$��v�Ukg�!�7�l����n��cs���g��9K+$�����Z���@F�����}c�����\_P5&o�g׃�מ.�O0�B%��l=�Y��Y�}��/Hݤ���6W������5��� ��5�}��wv"u����$1���J�Y��x��嬽,,�'�®~8��3E��j���{6�����xݻOH0�U����h�m�hjv���Jt��J��J����ĢB?-��q��A@��:i���3ke�ͽ��%���2Bq�pj�*2O9�QJ��@��!����f;@�֞��̮$���d7�Ӵ�\UZq��$����.�PP��_+,h0�SH��8Mq[TG"��l� ���}�nvW�5�������=�8���($���[�3��\4#�}e���Vf�f\�MR�{qx@�Hb6M��
kK��E���Bbg������h0�MŬ'W�N�'f l�C����y7�(�ÇW�)�5&��X��(�Y[�l� ��f��脲�L����Z~~\�}����m#���73ܼ�� �z6����.`����zC��;�4"��"�@�S�U�h����T���2�aJ3�hX�D|����bWh�I�;�V��-�J
���p�Y8K�ŏ��[��>h	"�{&(�͆JD I�6�[|��]��C6]I�h�[�y�"�J��������]b���o,=��d�ֻ�Nm1�u�n�9���mv��W�T��Ϸ��~�5_�7)���X��!ښ	@��a����J�N������u7L�v�s!Cy<E���QƮ!��֪�|�׬�/6�2Z�J�<�E�i��	�)��d ��i��^��LIj�>��AD7:�ۣ�o��M�p+G.��>����P	ShrЛ�J0�[j���ʢ]~���ZMa��A
�=���A3�E��F�S��yS3��*z5�K��������^�e��7:��N���:�J?L���f$m��a!�.z1����G��{�X��r�=�N�t���	~�ޓ9d��;:E�;������WJ�h������:0�����Z�]�`���Q��^�m��yr�1��&L9���.K�Бu73A`c��'�
�\�d��AE�>M@���2i^5tʜS���+t���w�R?2�&��2h�����N"na�xEd7�����bH"�'s��.2K*�2'��������[~+��׋ًk�#�\I=�����wj}b���azv���A)�Z���ď��}������Ȥ���U������Lkٳ�L���.}L���%�E�c{��}qI?�?>2���"�TG��Ql4/�0���ԅcz'hesMrQ�j�9G ~��-Ҷ��<ψ�xc"�7���-���LK+|����~У��Tg�� ��_�ȕ��ֶoR�n�OдŚhy)�h���i�%xd�L<cs����G7NsTf�r��	�r�H�7��(��h�unbHly3:��&��^g����F]R;eP�1�Ƅ�ݞ�@<�s�p�o�ȫ��*a�~/�������r����2U2�I � U�C=�*�X%�����p{,\�4
6淍w����k��a�6D���pU�( �������h��Jn�1u��}�"Q�����YAd��P �������{/�/�0���no���ޘ���6�2��9���ɧFV�����=]����~��cS��&EP�z�"a$@�{�E1(/%�N��6)�<8�e�k��=���Bï�}A��8��}0����ڪ��E����]��԰v�����9�PbE�ڵ����}�.jL:�ςu���Å_�=�q�@m�^���g�m`�-�qS�k��:�D v����`�T?G:;����sDn�(3�� 2(2i4{n���,�nL���^�^&%����O�a�1plE�֤�wޗ��	�g&-��t!U������_���"Qn4���O�U�!�,�-��T���s�ug&�en�vCR���I�0(�}A;��"/�#���{��%n�������!�Ud0������t�B@��f�����<�F��Y��%Gn����?ŀ�$畣aӄ�W���ȇ���������K3����}�ĸ���M����̍��\oB�cn�겾P�e���|���<͂8�	 ����UON��\h���$���(Y;������Ʀ^+ҫ�J������<�Q��Z��,5"�]�萼X"-�ދ|컼��f@Y|��H�i���<�x�wy�끑@�&t��q�-ټ�~6�[�O3���<V��	 �K۪�W�/��_�'�O�K��A�|�ė���qe�A����Q��"��"���=\v�q�a�FI�t��S��g�!(H�|C������+��d]����4-�9m5������Vq�s�Ʌ�1�l�?�{G��Bj0M(�hh{[���� �5W3Pӓ�Y~��"1��j\%��.=��1%��.� �ղN�5���2NK>BdxS�=&��A�(L�z,u��gb�n)!Y"4��S��<������
 ��IoZ�Ҍ;�Σ݆��r�m�ΔP����T��m'�����D|���lDj��R3���k�j2��$����ro�ĎS��pO�i������2?���\������L���Q8��vt��i-��i��e92j�;�0h{�攍����1
��L��O�p�pA�����J�}�^������ŉ��.��4\��y"j��Htw]����fr�_����Ї�N$M��ܦh�T��\�ۣ��nպ�q�'F�����d#9w��t^:�䇖�$y�mq�8S���z��eq�ɟ����@�م��+��dM�"��Չ$P���{Zh�#V����p����K�7 ;��FKq�u-����d@;&�Z��;W�$@]v�!\g�����Ҭ���E��l�vazMJ0ix�vl�U2����3�H�گGL������r��.u�z��֙d���,�` θxg��e׿����	|�ϧz�pĝ�-�GU�a� ���
萡3 3;�1�i.Rt�Vt��-���HM�'�*aT�!�^B�u��G#���?��ꮛn��j�'f�G?_����m$���$�k���6��"R��xzRg�*�L�s*�߫�Y:�O:�����:�:����`���N�	��~m����/�=�U"��J�"a9���\{�����\كA���
.{��s<�����/r�W���	�g�:�8X�Ӵn����N����Q'L���}*I���)��Դ�'6b���Lvxy��-B	Ǭ��16a6f��G��>,ɎL��BG��u�q�<J�s�A�R߁$��W�����s���Ҏ7�VH��`��D���,��+�^��M��p$vFTuo{�� ��h[��E�]�k�g�W��(�h�z,�V��~�>��p�K�z/0��*XV����1b��xR�[/�,�x��4��%��b��px�JL���Aڑ9HJ�k5�Rq���偓=�п?��%~Fڰk!֮�N� i�2o&��pm��v#L���Ո^�,t��\��R�#�_h�_��d�{�I�{�1���i� �r�qp��UU�q7�Hޫ�����T�_�NYH�Պ�9Ln�`�0�Z)�uz� �UTS��(�^�4§&���v@S�uI����[+ �����M���ݘ#�u���M� ��:��Qx3��st�7cy4�um�4
�-�$M�\�`m���Xl�vi�mnG��/ �Q$P����{�|$W�&����ߥ��8���Y�>���G�
�K�n h�
o�g�f�Q�Lw$�6m�=��ҏ�(?�m�]��q��g��~D��5��)���UN�������c�YX��|��*�w���CAXF��<s0eLڦ8���_�K���2c'ROF�<�� ��j��Ρ��`��)���ty,�ؙ�:�N����)���H��{� ��O`����FVr����\,���s��!a�|
���5�@'��T�{"�I���
�P��H���?���(�����c�Cɦ�Ȏ�Kd�ܖꢠ�-�A�F�<���Gpd{U�
i�?�H���9�&߳Ⱥ�PJb3,HB������v��d�V��}eiW(��!�)���6;�	Mo���$Ĕ E�=篆Y��[3:sg?�a�¯�̱�D��sJ܎��헋d�f��F���A�)�2ё&vg�|o��Sԩ�M$Z�Ў�N�X���I��X��.��3�)WO��b�^�"�4�U�� ��Z�t3�$w��@��&�,r)�l��{��b����A�{��n�A!`QQm${0�ݘ7�O���%��Â��*�5�C&�'/xP�z���-!�مI�G�����$yUpA.��4I_�Y�p��2��v��i�T��USZ���ad�P0���/�(R��_Z��Rm��d�5Q�I��o�љ��t��80�.]�w�� �d��1Dd��3�\s�IT!� �y�zBMG� ��/?L%��`7���hʧ�0u��GjS�����12Y6�äO�*���SW-&�w�&j;�����f�JB
ψ'Z_�a�~��y��κJ��VA� >�ON��_�^��:��� �1���k��1E.a6I7�}���d�M�]��k�J����Y��"��R@=$�9��l�^-���l�Õ�����dJ�a�(k�\����}m���:�$b�W��@itaG�S�(��&��r����CX�����qy����>'Sb�JGf1��|z��w7���%�G�^��	�s�p*q�A5h�=�H@np~ �i�l�x1��H���T�Y~��nPT�?�s�gb��'�`�������T�kU|h����@�R	2m c��r��4oJ6�D!�We]�W/]7��#�8���8ғ��_z-}�AY�mm����W@��^�k��Ouw�\������)�sq�����| xI�̿-�Ț!҆y�݀��.a�k�[tK=�����2���|2eE���jak_�*�ՎM�����~+nz���!R	����X���x�I*37wTUZm	���:F1���q�_���e���Ԥ^��|	"�un�a6	��ǀK�Q�K�M<��ї ��v�����e�{��G䮀S�d�������Wv��p�U�l��KMl5�v�赬Id�(z_��A'�� 
K߉������tKx�(\��	��.�(���P�yf%mᘯ���=�eP��&�v�h�ƠO�#oimOfu�j(W�k�_\8��醖 2+��Y�^�6���ď���OI<s�L���PɘYF�{_���o=%���E gG;u����8}�B��$8���H9��TL��?���w"Ի�N��s�B�Q��l&�qn�~�FL����&}�~�z��`w���p�U�R����5a*K�	��QL=���X�Y2
J�:f�����?�i!�k�a��.�O* �މ;��l�K%��+?� ߳�*��EE���
�M���"Jd��eZA���a�=��'�8W"��C̠�S�>;��tF�_�`��Dn�M�(Q�U���Iz`�u����`=�W4f�5��3����t4圖5@w��U�oq���i�D{@7{T�����ŮF9	z���Tʋ-P�&�f�@�p���>(�8i�^��O<� �	ϩ���4Pz5R�;�������iyz/r�4�x�n�Xd�Cq�T�V���1*��ƍ��6�1#������ts���`�(��qs<U�F�_�L�I
�����=/mz���~`�.7@�O$�M��0Z�h\��/$F�W?$�Dd�&w�uɟ%��f�qix�*��s�D�R��h���W߼�h�����K�
Zp�WGo����m��_,��k4�̘�0�f5���?��ʹҵ�rj�%�-��g��ۋ��'�N
�No�0S
�[�"��(5".� �h�|{<	z�wqs��^�	=tgmm�yiS+p\,���A`Ӵ���fg)���AV���Yd�Edc���,��O��ّ��=<�0��1:�T~��3�����(ĳ�3�0�'��������X��g�V�s)�gU��6��0�'�}Qd��e�}�x�Kv�;���G�jĻÓ�6��a���v��?�'E������$��`�uB#;�VFM�e��E��g\��,Q��$m��t}
�n%,5�a_��p���1K�
���Eo@�q�WA�1����B�tP'�x����`�Z)�gɝ��l�h���1'��V@p<uz�cT�]�|�������&�n���[�%�ֿ�RմPL��N� �'^�i�lf�����Np�ƎZ2�L���z�=VMŀ�9��4͂;S~����Y���!�͎�䃫�	yt1�"�B�T\�kW����q��+�|n�r��^��\��#�I|�l\�:.E?7X�*�F���Ƥd'е�[�ƽS��7��M}�y��H��S���<F�{]A�5ȑ'\�v�˩���a�*f=�j�N.� ��i���P��4��: �vU�%HfPl�R�5U�b���P�4oc��[ �g��a/����!���H�a+!�q	��O`8E�@��*�[���x��ਓ)X�4����+� j���N*s��b0������KN}�
��	(!V�;T0U���{�;���T�&����v��0���yW�[�ؕ��J��@$�d+�;��Ml�2��H ����]�qzl�ڍ����v�-O�QѨ���O7,sf�����;F�,�
~=mbi������Ș�fv�W!G�ߏE��뉓�uh|w�p�8��8��]�2��i�S!u������!Uә�g�
��#���PmH|�q xv"_L�Ɛ �i��]n�ٳ �H!�- �ȍ{M;po�ć�m��H%H�>��k�aw���t��0��?�ô��w,��z��Hg���&w&�w�쪠�X�"�!'%�:媨��gK��e%�8jV �#�,dy�@��%��m�{A�2��%��}�ڴ|@O�a�t���b~[��kzlUKa��M3{�Ew\�X�H��滛XG�O`B���F�p=��=h�J�y�<@|g�S��� ���d۹�b{\`]1�(�E��E]
7Vz�˱�`"��p�R�Xӛx���*�։G���7��j{��Ͻ��݊&��M�p�P���K!s)D�2�~)n*���B�(�tЕ$�☎1���}��{mq?߿�����Y{�z?���<{���J�q��
$��1��{�ا3��c���p٭0�-"��Ŝ<nd�*�
���n&��â���һ�q�J'I�D��[��r�+���<+�2���y�q�,��IK9�}v0;H�j�x/���ke���a<�@T�ǀ4t����H���Dl�ytA�F����i��K�_���n���
��v��<��<w�f�	�K-��c^�:3s�e>O�-J��@}���#僀�"Yݫ�W��i}#�,]�w#y���CO cU��l)�=/"����Z#�KRh��=nS#�Kg���Hg�n�����.JA�|ow`F��)��X�$a�%������Y��Lqe������a�T;�7���+����s��}�� LC���x��Tpj���)ɸ.L �Dc篽��b(�9JѶ�l�,J@�`���d�3vx��XW�0�����6�)��?�ꝱ�d�e�D�in�X^W�e��.p�z��Y>nzs ZM6�3��(8-Hϭ���-�˗�^��ܞ��$���Ci�zLa���Gk�����6ؔ�p��:m9*R_�ÿ]4G���$��mH͌۞����E�����Od�:�݄BI��*~r��[�B��Uc��?��!���ͷ�㸻^{"-�{��y��=7]��vM�l�������H�5��B�&�i�{��+}���'͆ߖ���X�Q^u���wv�䀯>Gm�l�.�������	�b��
�D'����:�3�[��`!����6�BU�n��b��B2 �!&I�I�T5�����М�?;~F�.}�ߥ�]��ťKr���-Ǜm����O�Q��t��7�����|�.Aݟ�X�<M:6�����j�3����F��+�+a&���5�d^=��~����~����~����~����_��px���2q�}z붡*�v��Nyz`�q/�R��'�TBJcz��nX.љ���e�BP���Mѧޭ����;]P_��Ks�nr5�r�T��!T�#��6U(\߾�\�;�r�o��S_Lԩ��_D�NX�>�~�#�F��1�+���W�e�.^��{}��tW��$�����i���E��7�s7R��M6���tä�Ͳ[��6{��:��ft�w��:)��me��O�ʋ3�Z�b٤�I�2���s	���!��]�	��L~�tdge�r4���}���|��ir��c���ϥi�!\�#������R�!{X�+KZ�-"��"|�O!Uo�NWN���+�5$�Vۧ��)�X������zݙP4�Ċ�՟���&z���I�����o�L
�N��6��1���뢻NyV��|�݌��\D�#i�����Â
�4��������7j�|#�`�(U�����TS�8��,+�	p����^��j��Mf:K�s�"*O��{�\�����,�lN.ڻ2�����17����U	3-��t�ͰuD��W!~q{T�b]�8}��t��8�Sy��y[p��;H��7�?ZڛHL}�{e�j:f:�a����c6`p!/ $�꤆lBf�\�b&՛�#I�.�N�h�+;얞a+$�۱�t7�������6�;�kxW��y*��
m��Vb�:_N�KԌ%���Va� ;�輀�y$YՖv��5���~9��q������&�g�>K�DJ����\y��F�<ƃ�w �|�r�����y��b)3<?G�� �H��K���y�Պ��Z��'@_�]����KcKB_a���-��Ѷ6»�]��0e���I_��d�l��q�lr>q��Y0��4�b@�f�m�Y������w0�.���f�,(��A5�z��jK�Js�؇2M|�m��H��Y�p�N&Q�������Dn�����[��z<��h���URr��J#�ave��6��u���S��V"�s9WR�隆�,���w)�J��nA�_�N�����͎��/���L��_1`�P�o�z�$x�JZ���#;_*����)�M^[��ۄQ��=��ApO���쭔�K9Cv�~#����=�1�BhJ�w��P��>�F�cv��)�Q�fD,�[�ˣw2賾=��8!�G�5q)k�J�d���:
���K3uw���gjD&�Y*��}��G����U.����ml�0nM���\$��_~Mz�M�o�z_�w-Z��Z�Wp�y��>�9����vY]�����W��sS�N�o2_P
�_*�]g� d��s��(���&,�qn~��a/��kZ'�J�{�N43	����l��n�o���'���φ�f!̓�m 7�X�±��ey���p8���Q��?��<({&T$���� �h�ؔx��b�d6F+�f����v��S�[r-��wa [�Of9�����wN5���vg��C�}h��i�����
?��;�I�6��S\y��
fǿ��$��٬\'[�,>e?@��ƣ?v������	i-����6�Prכ`����f�ݜ2'։���l�!�*
/d��'���ü�*����o4)�vQy�+C��)ߡ��TV!�yҊ#񊆖2��g=��̚��٥�	��N�mj�}S�� |�F� �G��n�_��0h6v7n� ��=4-?�\���������!�]K��Y|�hK��ڱXo��}oBr)5���ƪt�y6�&��et��!X�Bb�aB�?}�����~Ո����k�7^��t��ƲF��K�7Ȁ����fEF��ü0-�!��f�8.���GT��y�$U��Z�3����	�?'��4��q�P�2��̬�jtG�Q�f+c�gt8b���*H-�t���:�7���� נ!t���04��iĵL�b�s=!�@i���ŗ������>�/񆀝?,:p�l��49����Q�Ox`���;��MzR��HP�q~�����ּ��>n
d����š�N�1�v���V�2�ޱ1�`�(>[��Є��Npth��̈́X��8zTC���H���:��A�U��p����UR{�K֘�J���o���s���}��c�p���6r��b��3:�κ"cYO�W<�(�L��;��l���p��o����l�$��	W�\��l|�!ܩd?�pK����
�&=��P�-�� �>�+��Y����� hS�쀩�_�:�_�CrH�n����=��T_����Y�/ޛd��U�O�X9%�o�]f��j�*�ņBv�F�0�ԧ��R`�q�ޖ��`߲	�J(#
[�%�_�<����I�Y��g9�-�ߌ2Z�
BU1��hX��D��3�@δ�r�-�UK��ENX��0�Id���H=��4R�Md���k�z�>������->%��OX	7Z��˘
��jCH�խ��OG����d.bO�,⣢A+�v�9��������~���C%�����~-��D�T*�+��߸3f��K!�s�p��3�a8�d���mg�<�~H���Jan�R���B����f7�eL}8��k��8O $P�>Ռ�A��#sH���1N��'vK��ӣl��g(�Ω�Q�:�z�g�%6�@��'�^�_���Ϭڈ�M��~�
��߲��!��A�F������q��r�盆F�;�������(��ƒ���28��
~t�rĞ�Me�qE ��U�p�s��a)��jԓզe5¾ g�!�N�������_ٲ�݉:X3�?�a��V����5���l��.��.���c��7����a��������c�������-��; IFL�`L�Ӆ �[�]��jG��AL��C�������A��Sn�k�j��~ϐ��Hl'�����ֿ�{
�:�[j\g�fHDcfn�_�ڴr��|��yOihً���f^��&q��\B�J�~f������s�KV�e���:�>�$��i�_��j=Wr����s��Zr�g�U}�y��0�Ya$v��nw��F����Y2�Z$=!dyJ0��=Pk��p�d	����{|Ӛ�z��@A���~#,���EP���rR�=��N�E{�N��jH�N�;�LC��{b��^ӣ���~g� �)#���A����䐱C�G�EnN�?�n�q�2ع e E���*}�!�a`�;eņ4�	�Lj�2�_9rǸ>�y�XX���I�:�` P�[���grea
����!����s
�W	��Ѹke*�Ϭs�u_�7Q��������64#��Uշ�Dt-�p��M�ټ�@��\k��50j��
��l��1��c�ֹ]&�ES��x�.#w�
W<YQ{$�����Ƥg>�`��������ެ
O"2��|�%�fb��q�� �U�{���z�%t�j틬�0q����1s���9�aZ����ELT��A��:/�B�����A�k�b+���0���'(�)�
��B�-�ʡ�#�^/�'�c;ˬ�Z@����qc����?	Sߎ�f�# �b�0鏅��Ÿ�kZ��G�P��3���˙@f4���@�09�� <&�m��S�N4ƃ�+���}�V��Cd0Ea�$wVq%d���tD�ѳBH����)*�H��e_z�-s�`	F�=�9	��7[*)wx_�=:��������P5L��Ty\_�C`Y��dIQ�emn����Ä��0�/�/�
Ku�D��=�����1z{.
�Kt׃�㮳�vN[!,G�yˆ�*���oS|�j�\@�1�wY� M�g���qyM�7��j���K�\r�́�n'VY�1�@����������*n��Y�f�x���P~�%�$ż���DJ�/O�1�^�I�ǜk/{��-�ÜE��Gf:\�i��M�������؇��$���?�|�w*�Q9���v1\���S2�6�G@za�
h5~6����d+�K,�·��m�ue��Tr���>���c@^	�j���
H���^+N_�E���B["3�-�.t͜��s�-���̧������~�e�'�_�=��{�U��g��s��Ѷ�������Rm���^V5X��MwI~,���B"_�
���<�O���d��T��S5os��9�͹�|�ٌ!��	nS��Z�g͡r���L��s���>��1�? t�����JP��Yx�I�ؐ.�$�i�1|[�~N:�|R�̰�C�o𮼃��r����U�]����SԹaӲiI��0(Y�I���I�xM��k��AX��B�8w�:�P�!���m���&1�g�2������&��'���$N�q��4_�4��mH��b[k}���`�a ~vW��ML�ďmX��O>&�.M�rV���"?8-55��9�����Dg�o^XY��wL���j#�m�I��r��ei��e��$��P��%�i������t`�]9�!��>N1�����;�	@_#��Z�S��3����/%g�]�76~�mH֯J�ͨn�
�A)J�?���K;�.�/�+P�YseА}f�7~Iu�FF���sM���6��6���/��s_J%��*���JͰ(~7�����ݦ�KYA�ν���jfg�m�&�׿1��g��$���1������v���0vD�$9"��xPtp�T�Ю���R�(d e1�{ZE����&/@P�Шs�
g���5�G��3��j��VA��"Ĕ��7�����
��h��m]r��
���8{+}��Kǥq|�P>�5Q�j\�oxg���~)����H��$�*����L�?��<踫��2<.�2�HZ��Eȧ� c��oKOQ�����6���,snq��i��,6��LB@��5Z�`dh���oC�`B�����p�ar�6E�ۋW$���a�^��3s���ҜS�5��{d�CǾ�v�bq�f���e5�����b� �VW��\��3�������]�'���m����Dq�1�~X�3���� �Q�����%5u,��'��p�B'�\��ҥU1w)L��B+�2rL��'��z񷁻8Ƽ�S���4���tpaUe3 �|��~c�0!�����Xna���N�^d7�)��YߘɅ!��S��`��ШԿ�E>$�n�O���mGmM�4w���N2;�X����W+{64�8���䦲��-�r��� $���x�4�laH�FW�7b��'D���s�0��g����s��=��� н�6L��
��	 �:��r�%	�2��رA� �Y�:�Gg��x&�Q�<Q��vxX�ȿm|������H�FKZ�1S���N:A�8�H^�-G'�kDHaxivq�Bm��[)>��Z �2��t��G�nK��J-L�.�z�/�7g��s��B�S��,�W]�[^��.
-�t�ӵ��>ʨ��!)1%�;�o���!F��[wu�<�B�y��^K�X���J����P^#6��7H߃{���?�+���E�垫�]�,Ow��\���n��(�,�\P��n���}���s�sВ��/�ث�/䠙�G��+�"��$����oח���$�s��V�v:�$��x3|�v�3"��v��@GLj����:0p����S�w�lA��@i�y6q�1M.�$�|�a����x($�k[z�&d[ۃ9q��.�V��xw��v��E$��/NT[��V̀+ȝ͙�L,��ݦ�wbXS�'gf��rE�Ca�>��vbr��>��b�k�RV#��Dئ�Ѝ�ݪL���(X����6��Iջa���u�x�S���k�'�*C��3�3�T%��U�����'V������(��0�]��f����΀U��#`9<#zS;?W^�yP�QF���<kMG>�zV�]��nw��_.��z�����Q8�����X���}{�H� �1%�[{�p+��0�_NrSq���U8�.E�*L��]+�qJ�Ң-��#��;�JV��@S�%O�ʻm��k�)�$����"Ķ��$[U*Qm��U�Z��"tJB�H���c��Z�=���Hà�8���<�u#��~���~(�|�����),r�:�=%4�5�F~���"�Ũ���P�r�iq�[��`@Qőr�o��J� o����Ҥ���_�Wf$���*8�[Ė%MMК����m��?������9�M��'h��#���pfZ��%k�Vn�a�G}ʲ�3��"���z3�~~H6:Pv�Z0�3����H,�д�|�&�=}}T����!�A��kб´�%g���Uom�Z��W=Y�a��c[�xTR���V��w�~���fm�&�p�����n"�������@��2-�F���_O!���J�[��`�Mj/ �^�W�������=�	����v�oq!-G�ݗV7�9�h9T��y�9Uٵy�!L��L����#QV�,ceS�V�}�~$���]�z&
��R"V��gb���l~�3�hv;�z��5w�o�e�ҿ��1-�<'�?����t�ݪ,��*x���Q�Z���1�Kpjÿ`H漂�+eeW�#�rC��+�ĤYi� ���S$�=��W���;���
i�ϑH}6�E��>h$b�w^ۈ�gg<�PR�m)BKo��?9���1�-�9.��A���MQm��M��x:;��ib���ͳ$�R�	�X}��Ԕw�M���*�;�=�;��� �Њ�ڊ	[y{h �*w���i\	�(U�hX�&s��b�Yn��$�0�'U�,j�뿈��`�,2Im)��ƈ����&є{���%��5Y)����E� ц��Lɵ�!2$3����M�W�A�;�x�fG��#��8��^�e�/�~��~��&���r�1��+���T�ѭ#��mm�q�Fb-A�MDҢ��������9�ߙm4���"Ϻ��# ��Ru�E�0����O!�%5ǵ5���ZiV�*ň���Ji�/����Gz� �Q:��۷W�̈66'�������hZN�l8b�m#(�f���O� ��\0�����w���4qVۈZ�&�/Pl�6h�F�|��U`�'�&��h��Vs�U�������H�_�66����1&���D7�ma��8(��'Am����`�|��L`����ᜪZ�؈�m��֖I�d�r���!��`���u��WҐ����x�E��$R���p�4�$��dKl���m�\]jO�5��^Y�$%�!�?���3[�B�v�r�֪0ls�N˥r����Dp<����Fù`큒�F���+��8R�S�0W*,ah����-bN?�龥M��h욢��7j}�(���wv5�^1��$ x�PK�y�E����vX3�l������,�%� DY�;ąj��Gߢi��X�O�[Ғ�[�U��T�KX���5�x��s���wf&کh���-�^[�EY�ϟ���w��H��ȓe���=�|��
c8	��^[n���,�#�e�"�s�-1,L��;I�M��ͭ$���b"ZAQ�"ʤY���U�N�G����-h��3�F|�J�l�*��Iq�$!��4B�Z~�Vp���nƴ��
�z�N��UԨ�3��T�LHq��ʈjW i�GX�����$?�'�V���{�S r�C-;[���+3J-G���7����#�.F3\��c�6]��ӥU�"��C{�G�U�����ch損�׊��3������-[���0z�a<�=�x9C����"|�ȼ���]�n����)²d���$I�HbT՟\�칔Uo	A��̳<��0Aq"��D�o��~�5� \�Ÿ��Z��6T�����羆jp�旅��Iڴc܆���Ί�+�lfب�Mjm��DOz�n�6[���hmdI���=�֤�䌻+�3k�?��v��pr�����+=��k�،!ѓ�|��B�-� l�F���[���(\a5��n��^;�I�*1�,5�ܱ�/���2Ȇ(6�W��j�ˎ/���ҵ��:1�Ck������l�w6�s�g=Uϸ⡇gL��&&�f힮$��~�>����@9��J�D�H��������`M��*�+u�'߬�WX �%�3)=o�*"���'0�$�q̿��$���u����'}�!�����&��z���C���/��
�O?��?^�p��ɕ9r��S�8(*H�� ���|2Կ�}^���	�(Q�H;�R�BGZ�ù���hD,q��T1�S{�{�-h�=2�"j���F�J�t�ƿ�����Tv^���m�Quf1j�/>����YGN�}��zw�|�m_w�����@���q��I�qF ��'z���HǴp�"��H��O��B�1{�!�oX��`��k�C��v�8^Jpa��vs;�q�!󖄡�#����S�� �����!�, v�.�'�R�}Md���Lm$�F!'�Q ����j���
�z��2D�ȏ�n��Ӣ�m����ȩ�Jr��;;8��Mh�n@�%v����N�]��' ��9C���mb�q��o�t�h3v�=�.7K�?��5�U٬+G�O!y���P����2���V�!
��?�)fVQ�pÚL'
��}�x�6"��\�,��+!��9�+�|���Qe���X?m����Ϛ0�T�"��JGd��5�k���k�gD8�����{�$�3t4K�	����ؠ_��F��y '������_����3i�x����Rg$����{��oo��ˁ�˒��.�@����X���K��^��\�]V�=��ȫG��\Wj��_�k���RS#������H{�/X�"�i���a\��.$��|��0Kj �L���~�-�ЇLRY?=�X�}p�,� ���Gxwd��|a�$g��I���J٬��@�Gʦ���ė���Fi�5ZA�J��@��ܞ�Vȴ��VFL��Zy�6 9���}u�-���5߁����P5��T_%�;=���,y�?8R�Dc!w��1���~L�H�d\	�D6&-�K��zj����_ �,&�X{.��,�Ď@vZU�;�.�j��t��~��dᦁq"�m��_1u�4���Y�����/���n��h�ߓp�(~���w��v��rg�,��F�K4��#`����=4o'
��X^��c�eh��L�E��q(����UT��PVx��˶!�MsZ0�Z��n-� ���|��[�-i�B�2�3�����J���ڂQ���������l���2�~�$M`R�b�A�}z%%6�uv�����џ@�=8�1
Z-n-�Jm���m�+��NF_DKv��֬@HUk�`6�g�ԟ`���������2�aU�bU��ki�؄�$��3r;�x8!� 1�em��N>!3����0J!%s��uY�2������Y�n7X
�M�tw_�"�y<
���(k߲���+и+L=�3	U�ކ(KZ}U�����V��J�}�d�D\���U��= �>^��Ô�;e��!@:�\ukjm�I���v��d��7�Ģ%g��Pk������7�:͍@��_�p�����v�F����y�;:�^U
Y_�,��~��3b�~�T*��̒bt���U�@Ū@IT6ɜU�|��:)N����[������σ�V���F�:	�&h��V�K��=�2xP�x~h��'��dp��b��G�vr�z#�����SۅA�Bŗadא#����+���{b����rv;���'X�}��o{��E��7�$�"��Ɗ���q�׫��c�+^��|T#����(d��ѓQS,i�8��-��OJ`�����pW��ŮM�#MK��P�VX���s@�B�6䭵 ����_����|���[�$''d�-� G� -.����G� ���� �ʳ$24��_�Q�pX��c5�N��a�c5܈��_(�F�>n9ܤ�c�
����FǏ���Ӽ�^���}�|���y��[/_�29�O��$��o/�����m�Y���C7�$����9R�h��<+�>���~����4z�c�5#�ޑ�m?�Y����z��i6�ߴ$���-���3Xz��r�dd%,Ǉ����'���������vD���.�Z�hWuلg���0��o������Mq�Za]�?�yc9��k�rK��Mm�G���b	��l����\���l��l�U����7�Wr����(�SU�`��<r�y���/K����5�h�.�/ff��bĨڢ7�<���Q�@�6E����f�ȳK�"�0���f?�\���7]4����rX���JC�f��z�a|����9\� -�����R��9ߊ|]�M�l�v�D�C��N=NUB���<�DG�`Ǜ�s��H:z�2By���Q��҃�p~�+9�;3�[��ɢ���]=���I��-�x�8"1����o�ɛ�ؿ�~ɧ��%]�0�����ؚخ�_���%������P���PW���hƪ.iR!C�?mS����U��dئt�%�¦כ�c�	ǲ)��`�)�ft��&��UԤ���[�:&��8��p�	G�RR�NQ���.O� �ňİ	^�)��x�9�տ�7GȲ|=q��Σ{l�?ߋ�P?�~Zy����D�yW>�%S�߈3H0ݦy>�r�,qna���L��o���K���g�$ݘ_o�����Y86s3�W�̀�ǫ+�ON
@�o{��)^�D�/���;Z:~c<�[�\�3m�ݦ�����ً�r���Z�w\آ@��H�G��>́X�_p��a�X��羅󆖌`�l���ֱS_4f�ޮp�������'��j��i�F���y_{����1W��E}�%�r�5N�s������Ʃ��?��x�P?�~���C�t6��+��m궳��5�.�~5�є9SR��.ǌJ<�0��{۾��Ӕ�+�X��.G�>;��V4vT���+@�gL�*ϛ`��������7eC3U��=b����k���~��/	�_;�1,?1�(����6#�.U�v����W-N�X�V��k��xy�?5W��~s�~m�9����Ei��~�D�V�I�?��m��saf���(��#w�B�v�LK��|���8��UTL��k"�iރ��P�w�������T0�	�1��G�JFxb�)����o;�[}rd�ޢ�H��~�)2��/�?��i��Aq��W�١��C�{)c`��������ץ���������!�Y�ȯ�Oh{M�����*��n�8��'���xg�H_I�ȈP~�_[(�׮.G����ZǶs��Dψ.^Tp��S�U}ԭ�-k!\}��J����[ژFy>dn~��/�+�������p!�.��>n���ӓM�����h�O�W+�
z��M�~�em�d���f��ی���d+q�ɧ�[8ˇﻄ6K��P��7�p��i��l����F��6��ԕ���y��Ŏb����?:[~A�V�2#'?��W��k4ص��QZ���]�h�?��
>�ox>��l��-S�G%T}���ٰT��Ѱ��ی�=g����N�y�g��M�َ6�e'���ǰ�G����δz�J�zW��ޭ<����(|�6�-܌`ö�o������]�y��ٮ�@��M��,5͛�L�������/�]�������l��[#dC���O��Wg�P8��~G(�����Pq��[J#�|�c�if�ٲ���y6�U����Y�o���W�6��ƛ^ ��N�Ʊ���O��=˃
[�-�Gz�DU�'o��m�����q�f��횫6��w��!6������L��n[����0�җW�t8��B�?�l�6R>]�ӂk��`TNX���G���Tg[dr��*�?��y��xU���z���5�^�����_�dO������ĕLe��>̊x�yâH��t���=z�)�;��o�T9v����7.�Ai�~�)��\I�~�����|^=�=��l��yMZBG�kr&2��oz��A^�_�^�7r��z���װF�y�0?A�1Yɰ
�1y� �3�bv(8�I��d���\\�ͬe?����TF��a3���.�A��&1�
m�����P�U��/�ӉV�D�O����R�g�Lv��F5���=�i#�Ed��s�Ea \	�����[4��X��G���T��pБ2�)@�|�2��S$��6 ��wI���E�v����I�
!������n�����߃wX�Tt���U�-��]!�(��Ě5%�/�v�J)R�S��gPשQ��FA*|��!��(`9��=�.v�vh�xM�XoVx���34��-h̦����ǎ�	��4�~u춇ƌP�%d��������3{_n��t�M�ă(Y�e���x˗h�j���M`�o�h�ss͹>��PaR�)w������qN����Vg�4�Lt�(���s��=�y�{ �x��,\zlŹ�ٗXo!�T���k��F��jZ���,h�<_Y�Klz���P�|�o��GlU:{��-W���P�I���r;;�M���j/�"2����*eo��٥��(å�c�%;�h�5:�(Y�8�Ő�ښQ3{�~�����5�4	����I���a���Äw0���g�;�&��NƄ��=�z7�n����M�&�հ�>��T�O�-@r>}��{�ы�촡�w�5x�JcU»��ln8Ě_䀭4}���5<����=Ĕoa��w�ң�H����~u 巫�?Dw���P��e�%�����ONyﳕr�Q���YY�96�3��`��%je��OM��^j��<B���D����q��LS��5�5H3�n"�����F�*?�KU��l�P��eM�"y+������G~��</?em2peU?Mf�ZEs�8r<*�u�z����<�� p���h[(���ϟy�%+!�㢇|�����<)=����ss�&@�����E[��`W]�����ro�+��H9������a=U���(l����'.��۸9��e����o>yB0(t��L�����+���U�����*��␍�
/U�1�E{����h��wBygT�MU����@��~���bM:������z������c�a��Ѹ����n�T �\ny��Sh]���'��)z��n�F�s��8���^�eg���v
]1E�yd|n�m<2��T�f��������1HB;ꊐ(��#Ӝ������c�������N�-g��n췼9BN*�#?�7A��������R=hE3�C��:�ˑԊ�&˪@��p��/��0��htyJ�#�˹�v
i#8[�xs`ҍJpO�OD�A�r�aF��S�Q�X��ks����:�`a�Z-��G�;_J�!�|���R�vNi��rӄ�~l��L��4�$�5T	�ԅ�1��%��6pb}UF���Ȭ��������� x9 C����<�a����]�^-ݜjr'�Ǚ�w��9z@�@.>v1�4�,'��K��h�L�i@�\ S5�� ����p�i�6��@�E�]q�Y'���XrO����b�����I����./�8[o4�s���w��<�LG'�Q� �H�<��xPprQ��DJw�	>9��۹R!-;�$ h�l�ǿ�w̢qz�;dYJ�Û�������C}yHdʯ�6�/��/�|�w"�lC��u7M���^�!Q�o+�l���B�e�P?�ʺ"DS��x8)�$��mǳ@Ea ��
d8Ȳ���8e�� g���zrɂF�<U<ւ����D!��w|7��L��x=5D�^��F�m2�@ǂZ�6������}* ѕ�5u��_��}4\�����#Z5���F[��/�ʼ�ܽ`ȍ��FS1gl)ȝ�ʛ[@\e�[V�(ڠ��hZ�@�t��i��@&ai;yS�dd�� ��NY�(��к[�xW��c�s��3:��H���]���_{kV֌��"�~vf�%��Ȁ��ۻ���\�_�p�w��5;�t��^�����G�}�� u'�z
s3�h�?,M���)-�T��Yg�P���֝�E�`C�`8��"Ѷ	i8�;:�L�*�y�UtGKp������H�џ8�4.�x
+�B�Jo�<Ў��S��b�GK~h>)%�V��o�i���)�گ��"�,�Fғ<�~���hH눭�·$FD���
��QG@�gX��,�a2<����(��R���b�*��"�Fh��:Қi@��	E���ޗn(�K�v�kI�]2a�� @h��xz�EӷYq�������ݔK��.�~Z*���x��iqq��(�F�������d
o��.*Q��8��>�f�� <#���a䉥�֗Vx�LG��L����]����>ǻ�R+��˗�]$.��?�N,Y��r~{�^�5�zi��`\ݐ?k.�p˿!�����o.^v���9�,�^\�7�r��2�C��f���{�"R	�Er�C�^�������'A��9#�Ղ����E�P�d��� �c���5!��rs~���?�<��P	�s�Qj�(��o�g��l�j2�<�q�X�'Q�<�~h4��-_Dx��fad���(��[D5����X_�������}tr�k��Ú��\��0y��k8�S�s�`d�?����P7�Ե�7᪸ \����Q\�*��WPF��S
W�ъ��G%��8նk��o?B/�1�3�����V��_P��a�ek�J�j��j��a�y� �Ϛ�A&=�׏b�l��TJ�
��0�q[�q����-�w4ԯ��J,$ �z������"��c�Va�Dmb�ƾ���*n(�w��!�'�Ќ�z*����%/��2�G&["�;�0 �������G+�
T<�ǢD�_�Z��兠�Y�' �z#C�Aɒ{��i�T�
�
X���T���a F����ź�TWm�DLE0��ɶᇂX�ĉ�L��w�=C���햇�-�?HԔKb���E$�~;��r��i�GAG*��԰S�'��F+���	���q�\�Qa��a��4�2�;٩�d~F����n��/Ka�@rj��/����eX�5��"��y�S	C�N�Y�S��a�����U���F+����Z'�8#Y�cn������?����������Ř������d��R{U`^�{g�%�l\q�fM�7�v��Se�V�R�3d1��}H��
���S��T�$IÀ���<��-ȦG�)&E� �H�Sn=�Է���J�dŹ��8�Q���|���F-L�z��m聉r+&y}~������p�n��iL�@B�S5$g�˳4�����nxS\�_���.�s/�h&Ҝ�Zp��B�e��U�T���VU��`�=H���������g��|88�]w0�Z�����8"���jx�4L	e^Q8#�WɠFI����R�}�wJ���2-����!�.��a��x+o�����oE^ϋ�k\���Pha��*+��Ȇ��7%>E��wZ|`<)�쎮Ϙ��Br~�l���`���4L��+��+�0ɪx�]��#.c�{zZn �����퐃�4S�Q�\���=��U�(��:<:e����y��۠|Ex-�FIy˔K+��H)�t��Pi@�p�_N)�F�ބ��H��`;Q��Y�0*Y��,h���<a���ŕL���5)E�v}E�T�l+^���+�Р�7Tܹe�70�Il�bAĒ�&g}�}�K+j�j��#l,��069b�)*�>}��=����D�Q���u:�7|w��]�.����tk�N��K��hH�����wZy	�Lɶ��P��Vx��\�kڷ�+ɰ)dݧG�U\$-\l��n���$-^��j!�r�5W7�N�g���r'l���鳽���8.��`���\rp;�}�f�#������J.��/Q�����:_��ͻI$f��Y�Tx���*u?zl����f��X�Hd��wٌ��Al�Pr�A~+�ū
����k�}�.
8u
�"X��z�T}KS�^����fF��3|F��ɡ�/���2��p�O�V�`�w~�fK���o9�^���P*�e���|Z�kǅ#x���.ym�0��w� ��U;�0:BL�WӣrYG���w�bHQ�/��+�zNᳺ�
w&��G�	�l
ts�ۀ�����h��0w��$�4�)������VTcKS2[t�����r�>��i���U�i���=�x]�l
�L�殖��<�R���RA��/$�}`��`��uZ �9�"��Y7Ƽ{	�q�2ږM�G�|�!s$5�5�%`4�V05SbqG���l��:p��+�s���+X	��,����ϩ�fz�!�Q�_!g+@�(��J�Dn�w՜$)�j�z�	k�-4�tf�5� z�/ƚdp��t��(�;��HjfI�dx��"ڻ}�s�\�]>ұH˰
J�/V˓�Zt*��{16�i�6z3<����KZGJ����L6� �u`���Xr1���5d=�W�-38�>S�C�Y.�{��Z�`fJ�Wpq˒����A�%�P߷G7��+�{����lS]Ǌ_x�F�8��S=K&Roz������/M��btڸZ��xO�ȉ B�$�Ƕ�Y��S��W8i���`�_%Wmֽ����=Y�p����`���z�M<w��ڵyR�-P~9�*]�Ɉq���~�p�^�E:>�.dpy=¤�BpɊx!+o��6�X� �:���CLr���`��v�'�\��J�<a���B�r��7��F�4��k���=�P�[��8�����U#K�_�o{8$yS`��9�7�&?��֯.ld g�N��7�W�_����1P��]��o��L�#�E�'� ��KaK_G�m��s}U����@�I7:]~0�d[��F����{v(l2aS� ɿ0n�<�`��+��+���SY� �������銛����`�)�/6sS2<���"�27��6$����e���MY��Z$�½��V�b�{+�����@����7����үf۔|��>߸�L��7�"'���mn�f^��؂Ӣ��u[%�D�5E	�o��e�K�Q�p�i%���F��,�*E�oZ��N|&sd�!Mm�Z��z��sKj=�|�uV�NA�ixܴo��{�m��@
)���_��N��4[+ɣ�tΉ��l�mǫ7�����>L*|����ɉs��qy�S��$����B���K"%^�fg��r�X?��[t�H����g Q�}o퇕�j��/@�k��^O}����MтJ�{\�Q�o���50maٲE�������4`�ˍƵ�Ao#����|�>
l*�O�ў��$R�ӱ�Ì�cm��r�r~:���ϰY��Q˪��H�a_�kSX��h	��3;OښK�
�ڜ�����x��e��e�����L�����$Xr�T�Ȳ���	��l�G�^ �.��i�6�}+_j��K����:��g?�[_�g��e{c�9�:w�g�.O�S������o���N������i�_�Ry��<}]K��o5�ݗ���t8��.��g�	?G5v��Mߡ������jm�%n�7�u)��3CE}�a�f@�?ob��ף_�6 5g�]Q��B�O>>�w1S[�y�~���YT|'���V0�i2�����o#����8��vc`/���y��I��ଁ�HiM���>%OT��\b28�KεϦ5g�\�vJ_`�c�N	p�(|�y��&E�����I"jo,Xl�o���;��Y]#��b�����3erB�?3�Eȕ��2�N��;��������Ǳ����+pX)-��8�� }� �O١����Rx�&���W�3r"�������n����R�����m
���H���Q��T�]����>��@��L]�16��`��u����Ӻ���r:��r�<����#BsN���,f�2gwc�����޹�"x�1s��f ��JC����:�x��h�>��I)JJ}��D�v6n��T��;>>G���N7/�v滸o 2��i"~����K�{r7�
7���&������ty��-_�?���K�<�zr��{�}��L{Q3��o�����)E�N$�X�^|�*�t�H��S��u��[��� ���f�:�fb�T]~�i�� ��%��@�� ���V�f���t����08Ŏ�'Oo�?z�q�#pe�@���o����<c���C��%ܨ������u�0dt��R�V�>Nf��c��{/�A<�Pw%��p���2��w�I��?���U�{��D�S�W��T��=��{yg�������O�ڜ�I��z���.�	���������Y��>�^��+�Oy:b���� ���o��'��ss��jQ��#�"�9]o��nv	�F9E~�������^���	0'u��#
�7՚��A�T���/S�)����Dd1/oʁp��{+`�R���;NmkY���&K���T]wX��^4�QD�H�!(H� �h�TA� WiҋR��#(�A�4QP���U"�IH�}3��%��y��Μ���3�;�Ԭ�z`q�Ƿ�d�j�/��b�D]��|���ߠ�9*���rr&�|5�S��Ai��}Eeٮ�4s޴��íQ��ޑr]�"v�x��<�����U���+��g}�*�����uE��/ܾC�������P���<�Չ�09�2~��'fDDGA.�3B�jL%/ ���_�M�v\���C鼖���h�IB�I�x%luwV��e4"km�|ڙ3x�������\�����\k?O$(��#�t^ԭ�h�-��v�7��zo��|c7�A4��X�e<�x�6���A��鍇}��)�[#`)OD�QM���)�^�b��M/�����?�9���-�K1i����Φ$���!h2~�:4F�pw.>N��^X�o ��T�H�dp��(Ĭ���O�8�
�/� ����E�W$������J���bd���A�V�Iԕ� j�����O��+��W�b�����65C}�Цo_�%�u 0;$-y�������۹`KA'�d4X2܀I<G������E�� x���%܁_6�rf-.��;��{~%�~#�P�}�%dZ����Wz�{�����L�9P� 2?ɲpY�,�Y=!��o��:B4���rvMHFE!߸�K�����q�0�K��䉃�}ˮ���@�E�!hO��R�v��B|�İ�j%���ˣ�s�R�&��2��fv�Z���=������"�0K K���)r��0�������McR�&=�����O��)7��!~)>zѲ��xi���d�7%^�J����}=Xw��6��(x���@���r��Jh�ٍ<��rQ�N�(�NA 0□e�Zg�<�|DyS9��+4[o {%Τ�*S�߫΀�n��,�Ҭ���|=� ?�k��y�$��3� �����J�s�)��b�o<��fJ���9����!�
b���^	V���ܮKhڤ��v��Xzg����t�~���gt��rXO�[?�{|Ů�Ó�c��ϯSdM�[pS����֙��z��W	���s���@(�T��ڸ�C۠�	�e�0������D���DW!N�
@P{�E��X]��������,��b������E��_A������	�׳	{� ��Vπ��DJ�66�f���Ok�^��N�zǷ^I��q�y����&�����F+��� ˽�騙�q6�Ͽ�����s�2�&
[%&-ï�.(�����������T8w�zM�d�~�I�A��qưbjV�˶�OS��[/i��*���ɢ�K���Z|%�W0�-�
�/U�b$ҸI�c#2�-薶^���SG��h(-�������pU�h������e��<V�E�<u-���n�P��ҩ�k��haHx�S1D��8�rOǁa�v�<s�C'�>���>_�y!H�DCH@/��؈3�+�z�Տ�(�HuvK�<jT21��J�'X0�ݪ����,5�B���j��PB �(q�;SY%�f�������^���$Q�����ձ���\�)�'���jk(��t��t'l뗠��}vQ6V�zaݚ�C�eg ���P�
�Ż�՟-��n?�]���Yz�j�NT'��<n<��C�e^L$S�_����X$;u��J�ѷ��-��h�n�~���sHaIT�ț�U?�!����`<K�Rr�1�ff\ ��Iߠ#0G�?F���#���>]�;�t��.9����0%7�1���?��"�F��g�����-�n{��tp<�/�0���qm����!�R���rT.K@5�<m� H���+뱃	�9��W�,5?�ZH�$
]�k줷u`���_�W�l�Bse�Ԩ9�+�7Ⱥ�$�>JW�o��_�Ʉo���RwW�+�6wP�'C6���3>���m3���Jw~��������P���ԡ�3i	E/��d���s|6����U�w0g���Y��K�j�˄X̢���(;@r�Z��rWȢ�q6�� V��ʻ\;C�!H]UC�b�GB��ɵz�e��Mg8K�[������0f�s�����H�j��j�!������2�|Syʪ�g�\�Fi���Ct�]��lH-��E�FC����o)N�����Ы�U���ڥ3l3C_�xΕu�-u�}����*\��z�؟����4�v�t�2h($���U�Kg�Fw�Ja��T,v$�����B���6BCw#{���GGk>͆��n6N��Z��^�Q�� Z�6l�Vǐ��_��E�V\�]TQ�ݵ@�^f�C)�[��|E�5F2�-��M��X����y�ڦ:�����=o��C��0	?МJ��A��[�>�[e����#JD���P*S��]��A?��
r�~1�fae�1SR�oY�`t���B����԰�����I}=�ϸI���l��^��=^��.�0dL��ک�؃������N
��/��6�Gw2<��{P�!��ۻ��T&���N_(��s.�@�X���||:��Ma/"�i5���tt�y��JF������Yv�ث~��'�e$b�8NC��Y��z�	k�fS�W�%�d�Z���j�R7`�T�:٬�A�x(%(u*}{Ii��?����V�K�`�K9�@�W	z���1%/�����˩J���U����L
��-�pz��Ko��Y�����_����t+��W`gU �<Bl����̪u�?�'{��J��~� )�%<iV{��rS�L.uKd�<R�iٍPr��a �מJ{�zx��;�=��x��՚{�3��WKXm������R�0\Ѹdӗ���$2��)�o�Q:����C�7�H�@xv��>+3�#pG ���;_
g#g
�a�D�@k\�3��	�ǞI��/��������(���9lzY����Y1� �U����m=c��b��骻����Ep�=)$�:�?#��z'z8�,*�U���v�k(����X����s2�yz��v D���z�*�HK�rN@K��^[��ל��\���Lsb�u�w�)n��g���j���ʖ�Ѣ�*�qȄ��<�,�B�,�b�
5鷚��s�D� �d�j��1L�)�8KΪ(z�=�P>��UX*Lo�$sx�m���)�`�v3%���vY7�*�
c�r��]ggX�~���^�k$�l�{�tY<tI/�2Z�b�=��J�J��r
���~��(��qL�.�7%�o;!�*�v���(��L�OK�����D�h9��{Is"y+�� �H���~`��֣_A��]ٹ�u-*��V�nX���ʼfr�Nݦ�9�5Cr�u]Q�.�S�����Mx�[�Z��$�{-u3����@�bOU��c;ױ�kr�e���@7�����9+s��h����in�y@��L�P��X�F���mY��>h���g��*�Z���<%�Ώs�'άa켖���oJ�Նv ��}��K��r��;b@����2����}�;?g����F��iMݙԖc�����h��"��-N��ڮp�y�X�EI�e�DRR&	E͍͸w�L��������3Հ�=�Pָ��ꁤ����|��ٜa7nΎ�d�E���gI~H�(�����nw2\/(<DR��"tif�wݙq�P�z��GkQ�s�:
�Q�<��;��aeƵ�'q'z�1�E������H�
����,<bN�ː;
A��E�
�˯׵�e�Zv.�(��	H[�z�Թ{
�͡>!`e7L-�����kĐ��}���8P�$�ЊfG4R����~��Kc)غ�R��Ӭcy"�S�bzz��2�Y2\	�:A�s!n(��}�;y
�li���#$=-��6�6w��ؤ�|�W�wxlSmr�Ô[��]3�f_5qr=��g��,��|�l��	dL���L��:�!O��&7,���j�(��(�U�"^��Sz_+��|�p�u�0�;}��M�m>�[tlk��<�6!9>�ʣ����홯�t˓��������P��K�Z;CIj������'��w���\}�T�q�N~���ǳwF4��Pt����L�4mU�i-ď��^�_�Ѝ�zS�C$�����p���0�S7K�&�(/�x�N��l/A3[�_� mh\�-�����h�d�*����;3�& .�hi�	��j?�Y./ŔIr������|ܱ�e�5���_��3�����Q��T�f�eh
J������c7��@��&�HjBdTp��ՊR|�y3�'P�m�L�mO��;q��bn����Y~v��?�bʻ�V��T�w�t+q�lu���Ro���������&�h�z��d�o�iI��e��NS�'�謠�����v~S��m���ٍ���k�6dڡ��̉�H�c�i�ɵ�`�D�2��|���+�#�^�ve�2�M{����� z޶�jT�vY����tV��I�A���@���ho���YW������ �S�g��c/�8�j�5,�O����y�cPv�{���{>i�A��8�=v1�Jถ�80k�uM'ue#d�(87[Q�:힑��]l�������﵌�UY���p�p��]�C��:B���"=ߙV[�>@��Е_FTB	���w�&'Q��,컩��$��u-d��s1���Tu�M ��fW$����~��	jgG&���Qw2о���h����9�[�Z�ֶp��D�X�J*�1(������\�]{2����]eZ˜�{�ɲw��8iCnւGy��[)�ֱ}.�>p
23���-K�����` �=g�_Wn�	=�\(����)�M������w�Y�!�J�FM��/�&�k��N�1�PJm5�>�_{{n`�|N�
�}D�~�G�=mZ	#wP;sF]����ye����pd1j�u�N�5��w���=���6�2��%8�+�����&�8�I�3����!�3��!�x���IK�#.�IE�ڔ��O�?�}��ǩy��xJ�����F8���4��bN�~e�n&;W��Ƈ�o�� 3P�@�x�D�E�h�v�%:}ss�\��>�x�qG|�D�Fy�p� >��M2��c���]��"7��gͼ��Z�J(�a�r��K����w`�"�=Vm���n2M�!��aa��Y~�ѧ�NgM�ou��l�����:�p�$9���/��x��߭�s�M/pn�Z0�(���h�)�_4�`pj5E�R\��������A�Z��3R��k%~Z���m{qjâ�oƗ�LM�_MI�ˢ�\ ��Y��d _�\[Ϛ/�7�H�2|�[�^�������(��l�"��S���X4�,!!�u#�lnvc�znH)�LgzZ�0|�c�xjBM���� yU�מ��͵���vc��cC�4�C�[��/J��;�K�m$���z�ގ40"Ň�����y�;h�*�Rre;��k��%Ud��္����w�H�i3��mEb�|}���eQ��=H}ф7k6|w��W�i{�q�`���Q��p#&m�+�P�U��8�Z����9�J�UM���Z�M��Hv��)����4�c_1qy�=�M���I��nqw����Q��<�$%��q��ʙ���`�gغM����K���R������:��k��-�����qi%��K�W�;���f�w�xX�2 a����c�&눔��5y�,�B%�J�% ��n�CDt����!��O�O]Y�ܘh�c�7����#<�C���+ F��`]��i�Rmjʥ�0�t,����/�-e[�3���$�M��&h�.\�[�}��5o��_�>�$���p���0]\�3󏺱ՊU�6��S^R�ˉ�m�Կ�0���xi�������-F�9��'EJ�.�tI�� ����ulI.fm$_�T}���	�����@{�Xj=�L��j��; ۠K�!t1����� ~�RQ�b19(L�Τ�7'�<~��ĸ����XLE(�v��L�fP�F
�j�۹���#W/���P�A� �0��!��>qS]�gv�hz8�Q'��4NMX���;08Gk�pe~�����iiT\x��UB-}��[t��S2�B¾]�v��}�h�_f�mod�Y��,'JL� ��쳔��OJ
گ�O|��ږ��9�v�֫�y��i�c6I��{f�*�2�y����_3������'��"Õ�[�~����k���7�ӊ6��8H�3s���pé������ծ�s�鍛�)p�D�&��B��c�u��l�)jo_[�-�٨�Am{z���e4Q�$Ƌ�مOI�i�I�~bEߢ��c�[��Ԏ�%$��[�.ʁr��lZ��}ݟ�93F-Ye�Z�h���2Ӎ�1k�З�� \ZZ��/�C�&�i{��_�{���wK�jhSyX��� ͎�66�ʰ\>Y������N)����^TL�k�c��,��p�3^@v�`2ng�_��(��k�� aaHQKlb�J�2�*�6=mb¬��'�	N���򏿳�.^��3U=4�Y��ݱ�D
rc�m�r"7+�*+�vP�ؾ$��g�!��<��t'�c��mg��l7Pn?@�>���O���`rZ �B�&Lz�p�o9h���H0ifm���E�lw�YrKZ��Dŋ]{FԊg�`DϮ���S��tB=:�Wq�%M[j�q���s2���wG#0����\��$�������@��T׈�̆��|�<YP��a�Z�N� �z���r�l+z�,�|VJ��lQiز�~��O��-X���j
�! ��kfS�z��Ļ����<�ׇs�A;��v;[E(Yo����S���-������[)N�d����-�mn�KßoQJTN3d�2�샶K���q]�A%�����w��)���W:ھ�9�E�����3�h�Y�Ran7�������L=�ׄ�[�H�κ��Μ�g6�Tqī�r���K$>k�H�4�3M�j辩�*����>?A������f�W#����z��.������T��0-�B��ƧQ��2_�>�nWۙ��:v�	OOdR�w��6��~�̮�+�ŷ���5�P��~�K���`�7Q��j�ɑ�]w���6&��P��e�ۼ؎Y���-3��|6SR��;�P����'ބ��K9^%M�R�٬��>��؂���}���W(A%l�֜;+�掅k�t�Ǫ�.q��R7�������:�k���]����������t#�"Q�"tׯ�u����d��.O�����P��Z�`�ijP��wβ���m
WV�n�m9`�s�*B��T�\�V�/gsg�o �t�>�슮Ռ�s�H�_�#��N�������'��p�4�~�ěw�����~οʤ���w?���'���:�y�}u�_����O�n��.ި|&��Z!d��n��ʃ��+T�/�d�f\f\<d�>�|�Ju)it��z夾�-�&��SL���w���A;j���A��xv�a�[?�Ө��L��o�]���ڰ3�n$J*�����d��\��@���8q��Yv�oÃ���ݠ�Z�����Q�a)��>���;�T�������%���;��,����5;h�3�$im�U�V�B Gr�֥��H̹�3�������9�%���Le���ߎ���M��|N��:1Y>�y$C[�����o�у�2����$ILWS�����r<g���f��<��%��!ѐ-����$�[Rɸ�+y�����	��ߚ���t�@����w�P:9h
2�D-���`Mi�8	��ƿy�mO�(M���圻�}��/����s�F������D�!ӍM8�Q�d�`��l'���K�2�ވ��/"������UW�试�x
H�~��yg��f��G'�%%��Ng2쯁4����ҹ�9��!�*�#)�6�Q��B�t��_+���ߞLo��*(�B�O0R�au���=qФӺ(X���Ғ܏�蹀/��*����CV�K?��6j�����F���J@eS�=�S4"�%E�l�+5�b��8h��"ٜ��|����]��%��`$�)��6,���b9���;g���f�?�F8|6J��A'�u��#�Gs^*C��7!���a�뒔I�*�ʏ�U^l���n�ǝ0�t�k���UG�����~�ZG�ӆ�Y~]es��uڬ��L1!��PL��wL`��E�YЙ̼O�ב�����������/˳��0K��3%ph�>��,��ǿV�sΙ��A���V��{�A��# @�)�cl>?r�h5N��8Hm��a�ݏ�'@��Q�m�[���]Wy�#`l0��i��4��M��Mq�F 9z�Hj�j�NÈ��7����MN������9v�K�3m���(��Qg��9f�^G�˦�g�i/��I�Si�Q+����_����(.��k�2H�(����D�y����!����k0�tU�w�}���N%�bs4sÊw�d�˖nAb��+t^93� ���
�<f9ױɬSo��*��w����#
C�����9�����\���� _���j��ր�(��>�%%?��āy�dx�r�b5�HI���V�nʇ��߇lp�0�쟣q_���i��f�i ^T�g��ĝe�X�d���`�y隚�9X�	�����{�hi.O������I��cqb��0PA���°@j4Nr	4����ns�R��Nå�?��g�Y�����m�������\�9�m ��{͞2_EnoY��ra6�S�±uq����P�����d_%��,2�F0ϹL:[�&��Cۤ�/Oe�a�:��r�u��#t;��E��ﴁd�Z�uo�����xi�9X���2�W���!��*�UW�S�o5�B��� Ǻ�G����2 Z\�|`9)B��pd���� N~;��A,��_ י�̆��ll��F��r�y�������!�L�|/��&�vQ���8��.����hnT0ޙ�|����4�5���$sr(^�����o�K�U�BH� X�hin�'ꖧ�:��/�r�Iv��A��$l^�=��"Vt�r��SL\Y壥K]�[����O����s Y�I=ۘ~��[��C%��D�'��NTn���A{�	A�B�Fg�Y$�kˤ��|9k2�&�`qn���<�?���V�H'�����/
�s�'Hk�D��t�l¨�N���6�'�E^U������\M���޸�,k�P������BZEy�-�x��3���B��|�����(�t��*7�&p8(�v�hk<QV��?H�"U9O�3�"l�O��͘J.S�^�(R@(���=%[R����IvB���>�e�����˲tr���c�u�|�����=�������= ���~~L	9��l�� �?gn9�~c�h-y����(�g1븟O�6(�\��Cz��s;������ͩ���Ig�j��BP�&FL�O(���͓M�S`P���e��FSTp�o'�Q�/�5�s9���Y�Y&�)�:o,������aA����wQu����Z�{�t�0��j*{�*2�UQ˩l'�r�s(l�#��i�o,;v�^R-���N�H����y��/#����ED��`NC&o�t��K�y"3\{_���z`�`LJ� �����L���q͉�k�c
x0R� o|�,6�SP]�^��娷�Te��zY.@~�;[N�&�n�j{�D
��No�>b<��F���Hq�\�d�Lq�(�#�m�F6Z]�UU��?މ�a�:ߤ>�eA_���+u���?��A����X�8W��$eJ�dE�W,�lb��9�
���{�l��$oh�l.R��O{x���B`!\��f� y���֨����|G�ޞ�u���#���eWF���O�\�t����<]1L�U�(\[��~E�c�ȇ��-c�E�%����e7>�P�}X.�����\��%���s��T)P6M�V�7"2�B����>/�V��5�Z�W����q9<T��(|^�	_�;gj����YH6m �5����Lf9B�B���|�����,�#�<Y�o'��)����D�3�L��i���(�
����<�����}�>����/9�nb���k77h� ���Qr\���R�-N���©FLK�F��W�����e��1�͢���2H@��$3"��L��̣��x"�tY�e=n�U��T�a��
P3Z�?c���v�L�׀�A� ex��>����$�#��uP���e�{L�cCZ_zȍ�4e�=�A뇃���{��ĥ/�ġխ����0��9�a�,A��=�t�3�k�2��Ƭ8-ۯ@�乾ʫ�@���_�Bc,�{���Qwl�-�r���&q�&�u�Ɲ�K0D(���S�
6�����a1�	�Ɲd���U ��p]�X,�+Tl<Q�|0@o��]�g�29-*�9�)����Z�b. ����E�,lT��2$�v���-C^hS���O�L�Vޒ��q��PQ3ڌD��8KŇ� ���	_���A��T�v�,r��ic#z�vȏY�z;�-�K�~?�6X*���%�Na����ߒ��hsU�P�S\��
6���.³H���4�u����yXlzMV�:�	�t("wI�\����.>���Y�C(h��l�ޑ�H�
�(����7��Ӊ"��K���п�أJ�B��t�}��#7�*g�l��!o�z��P�S����xwJ�,��Z%������_sǪ����$�N�h14b�2qV
>��s#�����Q\�v�XpgD��Ж�}e�]��	nЭuL���Ll)��$�������6�����*�����m�e�����=�5cK��X,+��M�%)!�_���k�%45�;4=tl'�R;t�y~/6>Ȃ�����L�n��}��	:��h(z'�V��c�)�����3�!���q�^�#�1k�~ิ�d����bt�W�1���D+����wN_x��-�c:��$�@�Y?����H�1S�2�TKsπĨ	j�\��؏�"$ſu��F�6x`͖� ��[UU�G�����ȵ>��h�OoLqs� �r_��j�����]5(քa�;�$�S�����*��l+g��m�r-���	�fF�f�Zs�ɢ�C��x�f(yLw<|�_�J��G�����_���Ϡ�&�͸#�^Vmʯ�
��:Pw��a�+t���}|4��,��������(@�_Ӥ��lFt��3D�saI ���-d���U���F^~�ːՋ����(Mz�lW��!��0��:���������^���n����O՛��P���'�lp�%���NH�G7|�a��)a� "u)ZKne�]y����	����(qLN�����~6�u�I~Ui�G����PxBq:��d�6ZKE�9r]��d���ha�tv!y7X�`u�Įz�/��#iePR���+��/�ª�3���ud��\�.�i�>Ѓ�C~9�7:|`�	�/��@����;"h�p.gf�[�*q�A>e:�`��ї�5��N�-�_��l�<��Wu�*6�ax�`����c�a;����W�Z���g�6	�>�Ӥp7�d�:���2:G��ot�8�3,nx=�ڀ����@7����Dn9���� n;�	t�
9�w�h�g�T�'��8��x2^�sB��t�)z�Rԥ�?}a}���%(NŇ[�����i��y�T  �.�H	5W%´%��a�z�&��j1ɹ��TNt��}c!�p�.���:Q(S� /�2l�� ﮯ=��ܾ���AL嗶���S��,�0D�a�u�.4[ �N��ܯIQ���P�, �v��Ƅ�Y�����iԃ`v�"������,��Z������`	�p�8ؑ�m���
�I��}�����Z0.�>_-1W�.ۨ�����?�U��0>�N��2/ҝ��`	m���n���2�I�dx���k"�OZ�f�҃< �/,<�}[t��-@)z�e��*p�d���G�Ώ8l�e��z��� u��;_/�Uѣ�5��ew.�ܷmS�W�u�~u�Jp�<Yd������	��+�x����?�Q?F+�}w0yeb�q���s������.��Zp�,�ʖ�]�B��<d҉���=i�f>Z��M�杗1;M)0Fܠ�rr����Ih��+��W���;�0a�@k�s��v�~���(q!{tx��{�_"/�.���<����"Z��W��[z� r��u������⇊��ڒht<?S�����4������������KlE���� oS3#��E��Wâ�k��
@ւ;l7���<	 ^=��UfiFc>#%���э'����R��wu^(ȋ��)�����֗Z4m�JZ]��=�H �қ�>g�� �l�ڞ(���^/������>����N���$�����z����P����u�[����[txc�`�|CSN<�jE�咾���bt��T,Әw�����.��+
�6�G��Oy����?SO��V`�0k����{s	-�u�F�YP�8c�q�4��� WKޚ~llu���eBh�C#�W}�����������/�<���Og��1�U4|�yTel�����v�w�ț})�&�*�ox��@ű'���$ �h1���'=��;���G#���A��?W�t����W��`es��P�T(Ř�wc�$ Đ�`�C��aq����?	��<��U#6O	����z.������Ur�(�<
4�qZ�����@��[�ƥ�z묪q�ړ0@G#�GS�|�cSw�f�]�l���v� ���zP�]��MSSݿ�&��>��N��n����G8Nu�M,�e�Aڱ�N���ew�vpS�[� ��9�?1�她^ǥ�u�X��S�}VFj�	J�������K��s��j�+u?��/=/N��y�싍 �p;��"]��E;��p�dyu6*����QF����~�����bc�/X ���p��K<Â˥��`k"��Oo<�*�3�L)g��!aS�UU��#b�exu��瀨�{A.(�H���ܻ,�� �2����}ێ6�R�	('*��v:����Q,1�79�d�F]�{�= +���`ݯw`Ƨ��{�%�a�8S��
��'��T�gS�@WM��
�œ���.��G�z� �v���t�d������4=���u��,��evڣ�%��"�{ea�jQ���/�]���/��=�4��^��@'�R��2C]��b���6DI����P�~E��1)��r�h��a�*��<A:�[�lD���Zk�s�ౠa��}dk�[���D��	�7�0�����hϭt`72��]M'(�T���i���D�%�;JT�dqOr�Y�[+�	'�r��_��T���>G�(�~��PC���Pu_jG���'�l;��	���4\\%ܰp�]lA*%�n� H� .��B;���4��>x�0$�Z�k�+jKQq��J��������,�M>��tj?��HH�P�}X�ݻAj���&!�~*���P>����E]��{=��ț����s�|;�q����'�͍��Pz�����,�{�y��j���'�P�`�B	~����M*	��M|��x"�`]".n�n��?�H�ã[^r�z�i�~*F�B/U��U�#��h%�
1y�ׄ�T������D �_���Ǿ�0M�ͨ
�ڳ�}�~��-�9/W������^� ����Y����c1�ͫ�0ǣ��& �x�e��g<���Y�U�c���_����7��֝��an�j���ZGQ�����Z�[&��T�lR���f�¦Uk�M9��Ϸ��OR�����(B�Oۃ����7�%��S�7ٛ�jTF'�TSZb��<%��7�y���[i $�@p�5��c��%��n	�VJ^l��`�/��?rs�D�ǴD�I��
��<�r����z�~$����"����x��|Ʒ������-<���ƉP:�=1��^��4IсmU3��wV5;��z|��$�C^MI�D��w�4�yx�$���09H�rs�|ص`��n
��gnF�
o���� �O$�28���!�������3�] ܯ��n.A��2��2ӄj��E8���������V)�c��2T�%� iVM�7dK�kS��I_��,��($&cg?}"�N�CR�G"��?��1�#��~i����k=�m#'���� x~�#�k�H���H)T�� ��b����Ӄ��ā���:�.����@@�8�9�� �~9�B�K�,ov;�k����O�e�b��%�o���|V����@uf����S�s��	c���b�d�a��A߄q}��@F��7!ҷ�}����R_;����[��~P#��}(j���o�>Ãd�eޞ�9V�v�AS�i��#�e�����74�z�N0 :�����V��S(�g{�z�T���PClݼ�M[l�E9�3�X:�?5UX�]���<��I��Jh� �R
�> �s�������SPA�Z�9vͻ?���'�F!��1��A#>O��N����)�M��~X�]��7P1q!�A�,|+���{�fp3��(rU+���4Im�' ${�S�Dǰ�NFS��=u�:s�K�4i>pn�/Υ ��E�.����W�l���)M��@�4u]��y��?ב�Ù?2q������4Y��TU�ܿ���x��,���b
C/��9�\�L��tpx�!�w8�ݑfmo.�g���&���aO� N��y��#5/<�	i�GHڽ0*���q�%�L�	k�����geی�ay�4�T������$[��߾>x����f�2W�MJZ����Y�p���\���R��9lhj^�_b.|��kH�3�vz@k�?�W�Si'S�-������3�A� �8�6L�M�q|���p!�0a�:���h�#FU�00�(;X9>i��o@��V���b�u��Z�!�|$}��#�l�M����vK!'4q�S SX�3��I_��D}
��E�W\�)�n�h����=�\W�.̑�|��/�������:؟i��� /Uד~��z��X=�l�cW���,�ۯ�0|P}���x�sN��`[��ѵ�C�g�]��w�#�W������Ǹ]�8��y����^�:\�Ҙ����F�X��:5'�����z���4W��� � ������/Y���΀?{��Ĩ��4#8XS��_�k���2^}*��?��L/���e&4%�4�mì� g�*�ڃl\��(�^JP/��y���0�� �{���k����U�T��Eg=�6�o�i3k�"T0>��^?��o�?m)Ef�����((U�/L��i�w�(D(zI��7�	)�+���I��� j]�sW�MV������~c���GH+7��2�@S��0U�a����R��C��G��� �mh�{L����P�@n�#%�-i?{�Ԉ׷��H*m�@�������R�7���!>��}�Op����[r�;9���A��[��d�{�v&n�e_Z�A a4�pE߬�C��'��	t�w���Q�j5��ξ� ��x�yՖ��N5ނ9�?����������B�n�+��N��A����z0-��qROQ�5�*�1�?���?���A�7w�t�Jڟ�q��Qh���@�B[$d��7%BkoL�tA��vF긹,:'@9��f�0�3�}R(���,�鯽�ϋ���TV_;~d�q�z��t�$�j=ko.h�X�Dz��!�ɍ�;�/pC�?�l31�Ӂ��9��2�$���\lI+L؝�G5��G���Px5E)�����#���$-�Aj5��H7�����ܱ�Q
L#�k?���[ُￒ4�J�k@��6Ю'���S)��]�B�}@ZMӢC��b˩3�h
)웖}l�{��;5�yv5r��$M
x�~���&%�^00�م ��(�L�R%���xgi�ފ���m��Z̓�;i)'/%��,+�ݨ�)Ы 2�u@��wo�n0�I-�r�Z�� ����f}����~����H�A�ƶ�%��m�*�#���N �>�l�h�Tl�;AQ�B�ms<��r^IL�f���v�8
:�~�ۄ��������z?�`I"��"��M
���X�ݙ��A��2�mbD$T�wTT��3���b��	�fF/	S%���=H=L�7�tK�m4�޹N�(��@$�Ѕ�ſ��*�ȉ���y����v	���Z�_���N��4B�XJ�X��&�hZ۫e�ua9�#2ə����!�%�,����BH�b��ECjGt���|Ճ�)��m27�� �*!AB-��mz���^-��+����7q�C�C���zˁއ6�n�:Ԙ�=8��\+KK�A"u��9�qɚ��q|]n��2�=�`���c��~�MR�m��;�[��|q���,Pv�jN�Dڟ�ԽW�%�p1�cco��D�yev��9~�5�I�B�3Ld�"��}i-���8�y~�s[�|��v	4�<�]m簒���R�A��=7r��eZ��/��F�U V��'ʮ�?���-7�O	+µU�ڞ@a�3�N��llzn~wJ��m��z��-K���BD�w�?w���tr�1u���,R��À���Ԛ��Ȝ>oY����Ly�� ��&n[l�I%sڤ~��+u����o:@�i3�Y��a �.ͬdE��F9��%���^:��]kr;� �V���w��>��=~OC�7%�BG �a7  �gQ����023d\ϑ�[�q����֕{�պ�S^�:EJ6��/�2��sޮP�3~wF��L_�+(�y4S��@b���k�y��0 �\��[���Y��߶0�&�.���A�V�#�O��������� �8��]��v�l�����P�*���6�'R��6�٭�Q�ɴ6�H'�݀�A�����/G\�:���b���!{�u ���o����I!�dm2)���O K��!�*��A׈�CHo�v+)����&�( 
�Ŷ�/h������g/Oj�;�<9�V�,v����@�=�W�� wn��'&�_�.$%�X�K0T��ɿR��M?���WE7r��r��IG� � 1L~� ��M�\PW��r�D�Jf�1P%3Q��5���0M��΄�U��J�a�Ӓ��M`=��қ1v(�кe9�!i�^�J��[oy�&1���騖��߈at%�ϯ�!��c"J�5&�eT�!�������ހdF��p�3��ʪd�lu���<�п8I�q�����f�� �ӃR@'ld�F�^��'���J��y����f5 =������\�_8
���υ�I8�Vs�;v}U�6ټ�J�&�$�q��<�WL�Y�SF�c�o!���I�����J{ӿϕ�^<�@=�}0:�V�>��5fd2\��KC�1&�ˤ�]����I5Q1� %��$�.g/�-dc�E��nl�ar8�+N^?����7Y4"�!PCk�aN���o47�1^l��1�IWy	j(���V�=�@���m�H��{A�@=s ��j޿7���ӳWF��s����Ea=���t|��V�:^*c%�zd|�2K���M���\�U�&�R�����=�t��ÿ ���/��|��j�=!�g�'�\��o���g����f�߹)����j�~��a��85fh,L �-�D�L�F���iY�G�d�B����5�j��Vɤ�H����xř��0�#�[���gؓ_�Q@���$G}����1����=':��<�K����B�GB��5����2��Ltb4�ѣXRB�Ȉ��&���$G�R�4y�A����k��d�%#�gJ(���<)	���qu.�� �%�݂bW�U���䋓�3�Ž��Ѵ��f�}���B:g���ևwO�ݸ�4�5ğ	��Ls	+�����2	��������]���Ӫxr���ga�1r��D�~<��u��$f7�� E�'�������t7����%�Ϟ�$�){�`̡ct�=���>?h�1���?N #�b�� �]{�?��F`JpC=v*��HF�/��O����!eT�ͦ@Сtfh�2@�T��;
�Ӡ��q�T*~��'O����4��X������e��
��H�z��#�d[۾�MD�U c@��G�f�[\����D���C�O�<��8FS�ȂCj")����0ߤ7|ӓ@�x˼#O�6���͘/��k�����싫򋈑U�[b9�O�>�nm�2R��CU�t1am���W3�3��1��f����?��Ɔ�����n%�%@s2�!�!�vQ����2�`����$m��cv�`A��o�������(U�mT<��	�k6ɲ�Cm؋S��L0�4n�*Ɖw�32���Sw�:�s(ö�P�,Ʊ۔�*�CI�wz7eC�p�&�O�b���ݏ �vbg(.G��O�r��G�n�r�-��7]��x��J�q�����V���gGGa��1����%��^�u���y=������$�[t5p����V����/�ѷ�7��0���l<�u@�t���J����J ,rW��w��o��WMn�F�-�}��yaԹD�S6�k�m��0Hlsܞ�#h�(�M�sDW_�݄��`KO�!���"6��n���ytF����f�Ф�����Y�"�KQ��(?k-��kۇܨ�-�,v>�{ `����˶��U��%��>�Z���x{�����u9>r!1xNs�e���ev/��ǽ�^�K�X�C�9��۰��\�?��: ��k/���R"��H.����J��%( %]��"ݢ K�t*�%�,%� �t�7wC�_�s�=�s��wf(��s�7	���'9�vi�X����H�>�^�H������"1q~Y����yj;�|OFC��!H6�;�`�F|��]A��CbDB�Њ�,ӧ>w�Q�Ts�{u��]�ѺS��ܰ4Y�	��=�1��쏔���L�����c�yi��Yw�ƆR�@'���DP���a|i�~�-�i����1���6X�Y��hN�"R.��Nw≡��U$��oP��M��=ڍ]S�v�#n:WD�+EI�b^7t�Qü#	Ult�l��ԑ�F���c!�5mn����5�Ů�{3� J��������:�i�9��8��#�6̈�L�i�����@�>�Eu�}l`���R	���c��J�k!��aR�{� yB;D�7�	;5�sCͥ?0�ۅ�6�bRo�g��vUT��8��ؔ����r�&cI6@�_��O!���D]�f�
U]�(��f&�nSQ&�W-E����.}���c?�f�p��뭭wd�ˠ�]�%��#Ԇ���Z�Zq���~ƙ�E*�H�YЕ����q|L�߼���uJL��h��PxVK��v8��n�eu�1��:OqI�����a8����lG�i��Q�交5��\N�g6�~B�U,��C����Ǹ�!{�w�=2_��	n!�'sd�T�x��Cp$�*�*q$c�v����qj�� �^H@_mmKt�Z+�|փG~Ş�J��P#�?��qj\F ��̫�O vf�������F�����o��8�0���I ݰQp� D3�=I�W��z#@/ �_��C%��,Ф9\�&m�ՠ�	,�'k�W'�b~�}Pu�<�;0ʔ/���s�D ���t'�u)� =
�Ylm�pd��HB����N〛�W�������Uj�u�y�%����W�X���<&ۥ�VӲ]�;�+�&�Ʉ<�5�L'3g��l��B�Өmr�z&� ��CYmM	��z+�ۛH�yJ�+�����F�x}�J�l�����*w������x��ä������m9T��zik7��ÏA�r��_*A�i^ʪ4o��!�*"O� ֦��x�����1�� �rq3���cs�{r��(�Rq0�P�nlc���wb[�m����D��ʢ����mV�MSl�.�Y�Ì��=���o�ѪK�12���8�k� Z1�fT�|�QD:�m���;����"H6�[�g����`�Q��C��;b�������'�..���� �``��Dx�4�"�H�B�Խ7>ON���7B0vX�ۆ��� }0�Q�zB�ּӮ o[��2�j���)�Ü��q�W�G*��v0@km�MA�שּׁ(~d!�����{R�GI{��8�x�Iu���Z�Y� o6��d�w$�7I�3����/�ɌvMO��?�j�'��a��)�܌��['D�g@$�C��{�8�(��e�-�ݴ����~}Q�� }h����7D��еH"/S-%+$�t��ZL��ag?��p��X|���(k����U-��n5<�񿕌`�a�����RZ��(&�w@��n�ŕ����9P��:p��+9=r��L5K>c�bP���܀բ&/���NO���D\��ӎ��T�P���@�\��˱��I��u.#<[�vu�aܸY ���8!�7��;Z����`���jT�3��b?l]��酏-�������Pf� ��1�^C���c��l3D��2��Ԉ�c��c��f���?<�҉WRs�
�3�w�Cϭl������L',��ޓ�$�p�g�<jl�н��Yr�h�tk��W��RȍIz%���}1a;�?�M�񕥷�����"Nf�&�j�r���%����RWX��3if#�0��mr�?�|F�˥NIdo�μ�X]�u����Ҩڭ��V�f��ٜ��wh�N�1�[uӂ�Y���rE>��K!�2G�Gn��y�Z�]�BN���Fg�;�iEO܌�l��%�*��B�k��LFH���s�`��\�����Nm�ۚ����ZLh��(��'R�bKH�[C)ŭ��]�1hA��JE��6l��%���6�~���f&��dG�.�-���ծt�SO2Xte�$�Ͼ��������pnZwj��,3��e�rKwƻX���PFС����PG3���v(č��?A�k_��5�Ԭ+vtw���7$b}�WuD�}��$�@e�e�ᴔ�:`�bg𴔣X4���MEs�����tQ��>bzz�h&-��V>�@Z/Cd�!~���Z�(:��?�`,��fe�Ed��\=-��z�����l�~�;3:��W�Y�'��>p@92��z��w�Թ�ƚ� j�c�.��i,�`\���(�>�c��J���jT�
8�y �M}��2C�#��9O<C����׮�V��7d�ȡ�T�E[u�9F��ͪ�^���̚�cNL��{<o�$,/Zل��_�-Z>eƻ�J�v���K�m����v'jm$gznѪ�ad��.������뙘bg� Q���>7��gE�E�X���d��k`��ȪC�����YA�Ze-�Et���^?�����w߾��;"�G:�eH�^}�WC��T��3�Lw.t�����JX�w������)�k��F��H��������59�g��~g����T��j-��l~����V��s	~�SK0��9�SɎ�9v��~�G�-ۤ�3��������p��S���|c��$?kRS� FK�.����3�c:���)%Cg��!�ׂn�/C���������T��g�km�u?\�֝�~⸳7u�J��^J�����f��@u�xT�N�����JG�!(�_պ#��NZ��L{I��x�9�#g1�9�!�!��/���\#ߣ�L�:Y!c��F�>r�������=��2Ci-e6&J�$$o�B�l�_8 � ��B�r��?�Y#G��^�|��?��d�i��HIIq��J\�OR�v�<o��U�B���M����&�����%�\Ǜ,�M�B5��+�?v��}���� � UD,�"熜Q�P_��;u�Mգp��X���֐�^��7���R���VMs(��������2!��Uƹ������)<V��y5O]fEr��\�G	���_���Opp����O�f�3?��_+����.-�t�q]��>���`���t���k{{�#�E�d�]U-X��8�b���� ����?H� Z�b5���mJݐ��Rtߤ~��Ӎ�0����.f֧�93�'�	9O�(P]��ΫW��H���(���C��*���y���_U8��#�p�&�ApP{Ng]�`�FpYP���R��v�¹���"yɖ:*<�D�G�ѯ:���4�f��.��:�֝�W�AWz�ZZ�kj�Dɳ�<fh�,EFqX<��Mq<�N �������;�w `Y{�̅b=3��r�]#�%���lh�q	S0�H�.���N�P1�0��,p� �޳o�n��!1��-"�@X P'����!��ZY�Y2+�[�c��CXP�:4�oo�Կ����V{�<�Ŋ��xH�?��ݱ�[6zB:����"qL��r؇�u���W~x�:��T{�9�i����~����>ڷ�����\6���n��dV19��ܝ�\�i�}*H�w��@��cr�2�_\�=;s���<17Mi�O��AH'#��p�rJ���V���1�g"�E�gk�O@�jəו%�����A����<�`�*?:��y�_\���Ä�e���4��}��
�@ꗸ�Y�)(�|���R<;k�F�:�\{�;�ѷ�&ڑ�H�����&�/�<a<��fq��ZD��?m�2�R`S�gR묁DJm�����4�-�S�f�˪2-�
ģ�c�k���	�ڲ�N|m�%-(/s���#��t��A���u�n{�|�̬�}��)*r��x9#��}�2~���������Q�(E�m\��	�[���
����]^�rr�[��g��HgrhǏX�Z�-��������:7+D�G���.;H�%����i�0X���]��eof;�Z��G1���	���;�$v#�6�<�ר�1O���h�)R���j۩:�{�]:��2�f{�.�Be�	w�Q�jE	2RE���|�L����tI~��)PH~�C���Fr�k��C�wF��Q3�rɔ">t8�s6:l��S#<m�>�s`:X�g���z<s!G�~��>ԞƸ����>b��%-ܦ�"�#F6\M����Q�xNK���'���3b�^ِ�4O+���L�S)uR��{�f��߾����2*����n+!x7k 2��XfT� %B�ֻEGǜ2��?BM3D����su_���+3kE5)>�"�>�^�jQo䇯"�2��j��J����ME�]fa)��OL�$=%@i���O܀[�n�US�<(�O����ss���P�ʑ䈭@���d�k�s!�z6�T��rt@�N]�xAK�Z�?%o�8��P.t���8��.�Ãbm�E99�	%�։Ěҧ ~�f��� ��z��>��fg]��ڊ�����6�&M����-b�w���Ϛ�ৗ�ܰ<��Pe8̰Нuu��_�l=�0@�X�zQ���?�_U�������xV˔Z_�ԷZ���|����bh��
�u/;=�1��1i�d�oEG�Gq��وDP��1�s�*�A��b4 �[O��KC�bU@��C�r���J�����,=3.*C�;ѩ�F?�YV=������b4> �d�+�l<�8W=��&)��L��T��m��_���Ǧ�tl���3M��Ʈ�4���r���N�Z�6U`����TkscQHH�M���J/�j�'�C�Gs�|����9tς8/h�Xl�8-n��^�HA$J;�B�.so7�&p��"\���S?5�R��Yk�n�
�Y��TF�S�%����9Q3�t����>O��I�}��z8~�PG�u�O�4��x}O�&���?��$�Ԗ�+�Sw��\
�I��#�E^*'�u?�*��'#S����[�#��I�^x��1��]Z�o���g���5��~! `$���Y��a�X���F����Os'����^0s/I޴ALʼX`^�r�7��~����C�'q ��������C�hf�
K��B�Y���WkiZ�Qkk�Em��̩F�Wmb���g�	�ϣF[��,u8*�r�y��W�Kf�)<���lX��뵗����.Q4v��$~lƐ���<+ �kjT��b_\*�ï�F��%4��^<,���ri��Wޤ`�!���CYH��m��T
}�(���(�x[���,�-y0ax��ޮ�<Uh�H�pͳ�#��5��8YQ�H�=�8�r
�Ui���NВ�V�+��vCed����:�MhdE����b&ך��c=ru��S��������f��	"-Z��cB�ң���s+:��_�4d�t��'����"(_��*���c)4kя��m{h*�_���3]ݍW	�
4�7h¦hK	Oe�\j�V����D����e2�PJ�ʐ��b��TV�/�R�,�TS�+�]�ӑ�ם�D9ԧ
���)�Oň'⢪	���C�6�/��ɓ^]�Ma�.7d�6��۵����m��m�����O��d��TR���� 8��o԰r��k|�l��`�)��T�a��d��&%�G�%ȉd���u.M��gx�������ԏ�W���v����q���ü��$ �Z=�0�D�����[cx�\��y���U��h~5�?@��c�Ȋ�Fw��{��Us��g�X��s�w�i?u��/�q�-�%H~����پÃ8%��J��佟��V����	�>��:����`�M�N%���S�'��@��#��_>��o��X�}�X�n�&LRpK�B�ǯ
�(3���x�وje���z?�Ң��<{�g��z㙆\��������0H���w��^S��Ϫ<������e� .�����.f*R	���Y4�������c�;?Ғ
� �H�➨"��4�w1��
����3��Jghڗ�R�K��f�P��|��K`usF�υʭ��1�}Ø�����p��Z�<AD�Ǖ�Pp��a��Ԭ�V ��p�O�1p����|xv�:�V��c��4ØP���\i� z�������?@�ވݤ.ɶ;�n��V�g�<v�Kެx�i%,�9���M��z�Ӟ�m� ���b�8����qK�`H����O��[,��&�r����+g�Bk)|L2��A�� ��-�Bh��u��\��2?
L����B\�w3�z�/ +Ɵ�L7�f���g�Z���n����i��C_�ߩz�
n_ˤ}E�i����(
�~����:w��1���u����"��s��,�W��VA��@���	�z"HV:�a��Ɵ�vg�j �i��y��}�ZY��Ӏ[� �ǹ�H�ܐ���o׉'���To|U�?*}A<�҄2���1+U��⺮�N+���-|p�UEJc��$!w�yx_(a>�'��4-�+AMMl�t�'
j͢�|a4��jW�u�Mh�_`V�D6�gm.��!(�Z�̀���G�3�T+A��+닽�J9�ի��V<�'l�aB̀(R���	M�M��eW��A:����*�,��.%�ǂ:@�]P����t1^#E&t� uâ������f�\��M16׃3���'�:[��� �O��_B�5�)�����'i�CZ. ˿�cR��u=��p�-��^�
���Y) JG3��CQ�b�6�'�&+`�8b�*:e�ں����3��Ccm�s�.���A�E�(��@�p��糫���L��{�LHj��IZ��ι1�2g}'/�Ms�x�q�n����˲�<�8e�YW.��`�SQ�ȱ�&Kf�ĉ�ؼ_h��/_:�����[�Dm㒄����⃺ľ0�=���[��p^x�> �=:�j#-�1���H�j�oBG��/��� �	�M5	��6Uk���z_�����H�
�GT[!&Y����OŋM�s����1�Ĳ�}�Dj%CF���[~H<�y�U��>��T ��N�M�n�'�w50�a'���b���8��.Y��f$9�(N�F?�6��j
�6��ػ/|��5�����B����:i���|J�+�{؞�f� 3�G�RZ
�SW�tT�:vsC`�s�g��
�h�p��a�`sLa0k2b�uzP��N֝b���)`lg�zcQ�E�Z_��?S��
���M|���	�Ӱ�ee�����)zx�W�
T{o���E��W�.��v�>{2��ds�WA�_>�����k#}0�癣�Ԅ]s'K�c�s?��m!=��'��N<ާ�Q�����IEB��/�HV&ƦH���d���Rjx��-ýg�}D��������8�]9�)��u`w6MX1��j9M:��h�8I���qh��?\��r����Y+&n
�J~T��h���7J���~C#&LX�AB��\g�TTY�-��:XF9�j���.{h4�}E����ô e1�=�ύp**Y��ǵ���cH�J4.�0��c/�Y�mt]SK!ř�]]�0}�r;$k5gO9�o�Է/����e�@~t�Jݩ��F��mZ���z[?��j.��?)R+��}|�����q܇�$��k��_q"����@h�ҤU��-��4�ȯ�2(ZՔr/ߛB�=�^�SYE-�iR}C|U��=V�Ch��*��q\]�R�t(,T���5v͓�,?�e\��/��1���}wӝ��ƫ{)�)���Fd}22�^���|����bȔ+,��k�
��s�g�X~(ǵ<j�.z2�,�aEm�~��L?I��]3Ex��;����Ͼ;��!NL6��m�^37)7�	���������{ݴ��Jd����k6���^��%h�g��d��$��զ�W�����PF���/�R1Ec�t�#��73�qZi*4S1.��,��t�̝:\���� 4	FE"5�O��U�PD�oϋ�v�e5�À�5#�=�8u~q^n)E�il�W�d�Z��os�O.�U�c
�Ԥ2���[��"3$@��Jz#�A�s����o���WSnirArg�{�ʌK?��{Խ�����Tw�RX�p5?�ų�����&��Jf��K�{7l�%ngzy���c���3�ã�_�~?\�R��r���@��[=�[ ����n����@h.K����MѦ��Bsޮ������� ���;0Q�J��0-�,Յ�N�u���l� W�Ҧ�U��߬�1�*���i�W'�JM_�k�� {O��S�n��n
)���Ǆ�{�c�#b�ߎ�d)��>K-���J�U���p
Q�m.��gn����<��`c�$�2�"իn��,3�m,���d/�����^��JC}�Po�$摫P��0�ݮwkԠ��+c�?4����(�`*�D��޶zGA���T}�ȹ��7���-,r������!�z���ev�?��_�tCfʱ�{#����)�\�ʚ"��|4�d�A
<�stp�V�,3���עc��w��/`��
��,04Te�Ua��t8��奜j(�^�!>����SyP����<�j�w����p�u�=�q07~�;󓅣Ħ��ir{��c�Yk	@�|,�1���fUu�C�7i
���L��
�H�h�-��xdi��Z��
$�wW��S
�/9���Zw!��QJ�Xf�=�y�8mzA�}�F|VA`��~
�YНȮ`�O���G���(Q5��e���-k~�9�,����V�;Su��3J����3k�O籬6�\������������'|u����i�{؊¿�G~ &�X��;�r��`#9�����~���h����P���	�m�*�����8vs +���PMP~b�Yћ#�e��m�֣�����)Bw1 mgֲϯ\ L\?k�s^��݋Q�K�K��/��Y�ch�)x���~Z
nz���6��Tv+q�8;�B4�s�&P��/P���a�&����A0*
]���O��=$9[d�� )y]��$��^ib��g�YXU�㹝��[�y��m=w���\x�
��Qiu*3�,�%0�iu�{����E���z�g[?-Ƌ��e��{3|AzKK��j��u�%�w�5U�q�R' {��IXg��
�1�!Р|?1���r#���EE�qɭXS3�q�(�{��V�'��PoY�<�w���-A�p�A O�%��c�Ե�F_1��Ef�����[�Jg;$z�
�������Ӕ��m^ p�NSȠ>�Re�[�Hd�?_BLov'�s�ep�+�*�y������ƾ%��d����w�!4�gZCÈfw�Y
�Qi�}�F�A�d����i5F��0�PW�BN-hI�W�~�H��qm����x�Lva�tK�:kq6�@�H;����K��b�u��O����v��t��(K!�L"��t��6"�6�x�L�'���Z�ev56f�?Öc�L��)iZ��t������pFX��3[oD�N��s���~}!�E���ԍ�uq2[�6��o��(�$�� ��_���f��<��C�M�4j���P�ы���7�;�%���ｅ����r]5S�|�pI|�)�@�����_vՈ})V��_��^���xr5�S�<��uM�Bu����X�}!���;KE�:����ӧ��L?0�m4'#����"6��`p��7bFR���3�//ʔ�z���Re$ߓBH��U���40'�	ӔN��o������?������C+�ϥ����a�Rot�����s��{�����=���� 5�?D�B"�L5a��w�zocP�w�"�Ŗӛ\nV���79n�t/�u����S�RRқ��Tz9�����%�溬>J�i���;�R�cMN3�\ci^Y8~����F�L��}�X�Y�Ŋ�F���h^(M�?UJ<'��#�Ǹ�zmE�>A<����9G���B�N)J�L�v]�Z� F�-='�$�T��#�ǁ +t��h�����'�'������d��˲�{�ל�t�g�n��ޡ,�"����؇Ky����d��@���H����gU�5�����:���Co��1Y+���h�G1 F}3�KOQ�O�D��;�@k'y��0��7�#��^��~��%ibW���&t��3�x�J��	A˪z�oKwa���@��5*Z��,�c����No)6K(U/8�6Z��#FAô�I�$�Eh�_���M�~<3�G�0e^�{�3�)�;��R��G(%V~�i������*+W4�`%���Su))�� OH`��&v��d��E��U\6�}�Q�+���q��.����{�<��3�YD��%JR�Դ��ɱU6���4�c;lY�� W��Et�Z3��3���9S�Rg�'�:�Xd�e���zt�%�m�Q����DJ5*��������jc�bfs��<l�G�~�H bI�ʣ
�蒹s� |i�Gɚ��l��n�2��T���at��p)Z�9�:�.��z����4�<�3�b�n�����Ӷ-ýV<��|>;�w������X�����,��Y"7f*Rv�F(���FrV([Ϥp7V�Z&��㽩yj��'�Rɛ�ب5:�]��5k���	HR���e|@9|ߠtv��i!/�Z��0�Eq�^�8�m`ے+Hh\�*[3 �d��#��_�΄o#��߄�4t��nYOl	���%��o�f3~$5l�T�W��1�$�LĘ
!=@�D�'��D�ޠ����,�W��9��\�ߙ㹵u�ǰm��^^�)s�hcW�����P�a�h�纒:����̤x�{O=����gj��������D��xq���F�~kWR�J7J�9q��jm���;�Z�펯����W�6�S�^�[����2�������1BpM��A{S�����E�b4�H���t���8��'u�p�D`\e@d�!�z��a��|����d;�Y��]�Z�ץ.m,!>,9X�eS� �s�`:W{y�n@�!�b�ö,b����P�� 	8W�����C+Y����w�b儞�-K�y^���9������3�?�WN��TB�4���M:ԥj�AOu�YS�Qt&�#�Ѝ�^2]�����:��5m�]oa�zH#5�]���T �M~�xm����!�9�^���JXА8ԟ'����P| [%��!D�}=3�c�P��+ 6֋U���Q�G�(QǸ����p����?�SR�xybq`�#0f�z�z�8p�{$�o�:�����abJ��k��:���s�ˏ��"#�Q.�X5[�w�j����:�{�¯:) i�'�w4:�7��J�����_O�,�8���ϐx�p�+sw�t �;g���K�j��d��w)Sڳ���Q�Mɲ.fS��d�n���]�'xW͙l!�!˭s�^�be���C���F� ��)1��z�t��
*���w�xd��>��2�`����Q�[�����e�B�ٚ��2��R���L��z�N���,�?��m	�xn'��Y���<a�yެ���M&%G�<J�fX�s�9���-��������d��FVP�#�w`�]�8���D�@�(�hsx���F��#�����T���W���#Y�#���j��݀��;��نV�#��/�/~|����U�x��I����k�Z��;SL{��&̸1�T����C���k�kW�n��wĊ���;KP���N�N�Ϭz��P������1�c�U�f���e�C�*�a�N�Ä��{��M�lŏӆ��U
b�9�uT�;���*j�m��5���tğj�>�����do�[g:풚�Y�����8���p?<y�M���V�	Q�)�:e�U�o����~�>��e�=�5����� k�&� �$��)Ƀع�h�=�n� KN[>�t�����N�]�g7U��n�1br��gӠ�b�:�7�5)ۏ=�Z��)iW�o��^��x�"��Y���#7�;�LLtG"0�#�!�|��K!t�=^������U�o�5?hf�5�?�)���sJ�K秬QsNG:�[�0�l�(����֤����f�4׽����&t ��KmԺ���i�f-��N���G��RmY��?>`�og=}�?��f�Ӭm;��k�wm���!����{Kf2�'F�tF ��[{�j��r�|F!�W��İ��}���W����Ab��G��_��)�gq2yJ�a���hF[+`5��"��d���7ͳ9����1���8��-<>1�<R����EQ�>�,�����&L�u�ެU?,h�t� _ưI��\���l�uG]�w�?�2���m��y�b?f'-�;�&�Y��S���H���u-S��ͯ�������
��������ؒƶ���&]�($��n�~;���q�/����p��<�����'�2���|Z_�͟�0ףJ�{5��@{;�iK0��LF�-��qe�C�	��X�kΕ�U�`~�p�~�K#=�,����̫Sr�'jCJ��Ŝ"�8J�c�!p�'��w�����V%Rt��T��s�X�bTc;�N>k=�Β邉�ϯ��Ŭ�..0��c�%�)��s	�_�V�å��7Ƣ����~�Ӱ�\Px@�t�Q������+߲u�a^�N%=�dՠc7bnB���(?A�z��	�'']q-6��ϡ>)���'����N�*c|�z3J8:d�ޏ`~$!h��w����6V�J�\y�
,�i�`��a	�������h���؉��
,J�c�蜊-9�.{�I(�߱��ȐH=�ё�gx�|#�{H{�a����s9<��"���*���ɰV�SǼ3�g6��ΰ�/�w:0��.돴m^���7��<2�doG�p�'e��G#�;￪���t���0��K�Nd����w{]�B��|��F�wKD�.p��Y酵tX5u*�k5���R�n�]?d���r�E�Ku"��@�`FM�I�ꢸ#����p.aN�3��N���������᬴7Gƃ7Z{t��F�t%-I��q�X�6?@�Jn�yR��@p�@�OƙX����L�ܜ���1���K��G�Vt_�P�N��Ai�V��;��:��v��ۨ�7`�~p۔L���	���S-<�-*��#�2��-�aC�4��`�t)S��?�S���O�N��`MG�����|�zL=��'��40ZY0�z�F����0�ɧ��h�j7y���Z`r����VŻ�2|�%�D\C��<s��i(��U�eVV�L�׌���軓0y�åWu�Mz�ޔ���<������D'��Z�@Bk�Ƨ�<F1�`��;-�[i���A��v��֋AB@-�s}+=�,��W����#�����l���5���3'��ۋ��k����Z1g����R����fO#7� Y��!^���צ���<�W'w����>�x��W[�4cVz��2'����8�����z�3�b��J���;���3��n]3ջM��Y�{�x�t��w׹�W�3��#��t^WL{4�j�L��U1�)���/o��o�j��}^���å������e���`6-��ݵq7�DGv�;*uG�(x�'�NΗ3%y�e{�)���� ��H��(�O�ޠ�:��t�[�7�c|�@j]X+����X��3z���M�����L{AYs�� ���5Ͳވ�9�I�w|)�Q�pt�e�5�#,��S�"�����e%��!�'�aϪ���6�+�:�e��ȹBB˽��gt.+�q!9�B�q��4������ ~��>���2��	t��u����v�zQ%i�m�4ji$7~�9=���5cHNG|5]��n��i8ظ�~��Fܶu���L������paİV� ��g݃KJ��?L����w��O���Ӊ��m{�T�Dyh�J��&�6�x�6�L�-���$�����j)�h��ԚY�v���1�p=��~flIF����0~�)����,�!� ���w��LB'i�e+WW�)x��#o�N�MR���\��ˮ(�,�jם2ƺaԸ���+W<㸘ܼE6�l��n(���/-B�Y_y��m��H�Me�`�B�P� �|DCdj��_oj�F�y�_�?ڭ�=\��^6ɹ�V��ps��ߙ��G�7ĕ[ji+%��F�m/�.�Ǚ��A�I�������w�>j"_6�y��|Co�4����ޡSNi�l��u��ɑ�Vd<^��Չ}�7�B�Q׻�t��閨�{�k����'�Gbj�3�U�z��@�^%A���ʹ��=�o���T��u��|��&"^B�D9�r�G`��׶���ȍE&��M�Z�����y�fC
�G�����������GY�x�/����/�|>�"��8�����ۧ4��h������UW`h,��~�kHT�����E?n����@"R��;���F�����#���;8l���9(���E��c:��,ϯA�H���7?΄�s��ik��:�	b�T�?�:+���X#�O�h?�#��S�?(��S]lR��#��U
l)���t_F�8;��-����V\퓉cVA'�3nx�2�YڻU$RN�.�y���1�w�����o�s^<�q�h����7\N�a>T�2���g@��_\��D{��pl�J���ی��2Dc�^����h����d&�.95�-��\&�nBPƗk��l9�#�8�{\�a9�P"M�*��rh;'���F�[?%���{n?4�����O�8:�S�cM.s�f:j2P�ɍ�`��XX#������_i�����IC
Hi���iRW������pD�kd�qr����<��b���uʯ}��^�p��#m�l��3+?��Z�uY��a4;�� �>/�y�Kl����9u���H�Q��\r��8��}������_�C����f�:9�jJdE�S����v}{-/�+\}�^� ����\3k�8�x�L(F�~���8�F�8�}=1��)�����.�^O,�{S�:>�t�D9�l'ᙀ*�_9m�m��'�ue�Y3Jl��/�R��*�N�$l��å��!�,�*���c�
�%R��F��a�娾!E}C�7���-C6K+_Q	�me9L@��޽��1�y��0-f-?�����h�;��I���X��(w�/�N���[�w�V鍭XD���@3�l��D�c�)ok^̓ZZ+�R�o,�1�j�3M�-[;B:��4���Ү������s]ҷ �g�UT��
�Ź�����c����E����2z�~��K���Rk����|Oc*Чsi��B�,��4���ucM,��$��d@:{h���R��<dF��M���ڍ.��ϟ���ĊC倕X�nӿ��W	��,�^3}ű���@T:ڦ��-��y(J�f��(��r�o��Ϛ]��h�̧�*�5���S���W=��&¬�!z��n6�b��l�Z�hA��%
����kZ�����Ȕ��򯇆�����Bvڽ��6���A�3��l��33��*0�]����1�=��+�<����]/�k7ǩ�`��jq?L=��N
{�hJ̈́i��	Z94hÛ�Ie_&�bj�S������o^������>7<��@�\�B|���Rn;�Y&�eꎖ�B�l�����C٦�����g��ó�QE찅qҹI���\%�=E�PZ1M�6F�m�I�ei���膩pȅ���JH&��LY��yQ���D�E�t���n�	�K���X���%��3�<��
k��Ty����Z�%������ ie��>�}����0Ϙk�/|'z�;� (��rs���kx��;`�&��~R^�~j�'���Cd���K՝�����	G��_�h]�P{1�j�`EI�n��8,a�v3e�,��������-�
`}��%�	��]�F��L���!���(����hQ�џ��-�7S���b��Z�:�P�ǐث�t0:шa5<@�Ga㳦L�b�GgX5Kܿ�����ҩ ��bڗ[7N4 �����!w��U�l�ó�Ӊ@j��a�go�,ָ�t��W\�������8pz����wlC��F��l.ʅ���(���������0F��b~�3(n�N����w��5�.�O��Z�:ъ�A��-+NaS�����Oa\|}�锪�1�����(��g���h���8�D׬z֛$�F�?\�G&��k����l���\	9���5��%�J�{�}��n�`b 01�I�]���I��}��Ro�p)W�ʩ�� ў�L�mˉ%���'Uρ����n��jʉ���fs�L�)��Ys) �}d��`���Ֆ����p��7`���ӱ��Os[�Ŀ�?T�19s@l�+�9x��m�j�ԭp/I�W�
'̜II�g��1n]��l'�&?�;�΍��>T�@B.���)�3�x�7�c#�W�G��ƴ
W_ǧt'#���]�Qɔ����A+۱ڢ�9�S�ݫ9���U^qޒ�ڨW�*�ok���ҧ{s<�����ƭѭ������}f%3R�6�Z��8��ɭh�`41�ga���{�}�۫��׶
n0�q=�>�WS��m����<��t�~+���H��r\g=M F3�<;�����S{��*���h���,j}-��X�G��NPg+����	 �?Wry��X�4V�{'N�>��8�o�@�����9u���L0[�mkٌhQT;�"�Ct�QAi�9(�--�-����.�Vݨ�j2��(���MR�G�{�9m�"�II����������-�8�V�M�$j:˥���@!;�9p�М��k�(��w����-����
�a@&�Y����X�j7���<��H��,>c��������W2#U���-n+���ְ�;pV�)�AT�2
=���*(��x��?���ֻ��O��;Mາ�#> �J.r����7������^U�;Ԭ���BKIR�r��)��(	2�&{��Z���ל�J�M�k�7���i���C�)�K|t��I��/G91�X[GF*���7ڒ�1�M��H�@s�# �؀�{�|8������֫�[��ڥ�����3Z%o��ӧ������ǅ��w��ڏ7�{���e�#�YCV���'ʎ?��y$�h�����R8⁹�WpT�OSe]h��S�D��csx	u�gն��HE�Y�F]P��@H����Q��9pSd<��^�7�^�u
OUX���G�*+��N�����Q�No~:{�u��	-+����C�F��X5�e�,�P:$T�M�f�mh[$�{����
�~���X�;�=U�%�~}nj0b��X�>���[�4W�JUt���	��+�a�Vv%M+vת�D���[))53zYv�9�֨ �ݟg:lB�#�?9{�����S���K5=���뵊W��⡉����i��i�p���q���h�U-�{6�_����k��Wz�V��yZc��	�L����3�`l?|����ܤ��;�1v��鑝�u.ۚ�����\��B���a@V1��x	!�*F�L^4�A������Y�g�=)=�YJ �˗W}+�=�Zc����MmTC|3���G�NGjw�[5��M�b2�#��]�d�0��
���/�ߞ\p��>��[�%�w?�@�5xk~��U͕��l�g�b'���1��TQ�/X���V��&�E��9���U�ou��z�>�$�m���=���7��wm����t3�=�F.+ߎ��^��-�]�Qs�����'RxdJD �����9r|�쩡:�}�]!���a�lN(�!~$Vc�WR��ࡥQ��h�p�.� :��} t �!8]��[8hYɢ�#q��<���)���=�:/�`2���lʡ����lzм3P�Cx6V�� ����*��uK'���dU�6���iL]�T㑹hے�ے���?��;��=�7�E��`��HQz��RU�I7R�ҥwB�*��"5�&E"��@(�R�& ]J���&���w�=�q�';;3�2�]wY����b����p��������ikHh����Ms_Z�dxz٠+��A��@	��E%Z4	���V���ރ�7o�-��T7�d�o�ε���1ߞ��`�~� ��X��u`��(@@��@F�^r��^q8�(=5��n��E�hŬ���jbp�,K������Ί�ڔ�x�Lّy��$I���.�O?#WreV>�S����^�e�_P,Ӧ��ybn�1����9�X=Z�`S��^xv�N��dOq~�i�J�������D��:��E���;��	"fq�%_iR�X&T���Z��[�k�������DΩus�h�T-)(2�v'�L?lS1(<�/�^�y{���T��m�L?���e��>�)Q�w��Tc�I�"���o�Ϗ�X�&Z:S��-�d�,�&�.�����i��Sڠh�8c9�����@�j���,n�&����Y��F�_�E&��?^J;���}�aܩ0`0�����F �{(0(�D�ޘ���3iO	-c�OSS7���q��7���EMXA�)��FJ�ݨ�Z4�T��r³��Kk�mͣ���0�c��g�k��l��P��U[�	���?�"\H���Lp��|����o[��9���P����#��H��a��s}���m���F3V��<aۣ�2\��(Lz�+\?l�� ֚;w6��� Q�?o�S0�pF��J��k\�Yf�K~��T-�ջ���1û]�_���6ߛ��<���:Z�o��������j���N����z�������d��n�J���B[�(��_(��hI��A��z
��6>�8�)��6�2)R��(��e��Z�=���1f���Ğ�l_)���Y�1����v����M�8�����t�n�J��3�`�2��-]�Rж��U&Ƞ�5�yG9��v畝^GW�[�*�f^��������?����$�(S@��x�7����>PA�6N���wv��,�}�J�,�(!nB����@��]5�Pe��×�]���1�N� D%,�t��9���6�6�e}���u���N������(��ɨ/w7��E8|l3҄�˼���HNUc��/��ߏ��!$��k,������5u�Iq���"�2�F�(�D��c-7Kk����9	�����,�N������<'eNH�Rf�ը��?��xq���QEc��%��`�Z℩�}�?�9��Br�l7��=`%�}K��^�7�]���#⧩.������"�m[��O��3ox�s��}
R�@�J�D�C��	��*���#�Ԋ�à8/��`��f��������R��W�^8�o����x�g� ����ի��Rl8M,]W����f>���΢����k��)���@'�� �U,���>d��A��,�Y���
�+;�,����<���%����g�cT���8ͣ�/��d[�c��XR��_��k䪑��T�/�1�/լ6XՐ~3�E7�¢�����ru͓ϡ:[Z�%� ���	�SWp*:��C-�펵��j��ů��S³�MY�0�v���'�Tp0/ kJfw{�c Z��� �v��)���h�To�����*?A���4����5�M�EEw�o"�풵���T��,[2�.e�nJ9F��p���&��-��)�jPI����|�)��|�e-��'������hx�ّ�!"ɽ�O��G�C�mOuGѽ�$�i��*��)�Z���v���9)��}�Ȁ�1D�/{�4�17IU�2ń呰{}ǥ�#���)!5�k�� ��c_��yF`�[��?�����SQĪ�����r�)�}$C@Mxn�:�^i��U8<�������oE��ڪ��B8 ����/0��7PR]��h�j�Z
&j��|HN1f��������ס�k~�JIۨ�
�
��¾HA�L_p�rG�����S6<1���X�_�O���cI/��Z�r����V��G,V�Z���m�r�vFvl2�'�<ܜ<��o��P�%T��#a�lrv�M@o��R9%���O@?�����Y��}G|�Ai|I�����I��d��+v��Ɉ�a���V̰�/�����;z���A�{Ӡ��w�4����1��-$��A�ʭ�0��l�^�W��~�8+�`���n�4dZ���9ʠ��o����9H��G��J.��@���ז��5�Q��)���n�o�3�.l��I�"�YX��z�D�q}�2��ֶ�&2D���_��D��E6��q�[��z��N�fR�.�n��nܑ��,h@�A��Հ�t3o�ɲ�����;�.��Z�'
�,�=󉽈�I�y�]}�z����(���{kM���m�ֹ��'�у��ͩʫ�{�ȽO��\i���Ç)�r��v�V(��A�颿�m���������f�v��Oߴ?��t�]�,�_�ֈ�o2�;�Q�c�������6�z'Y ���[�*�r��olB��{�t��B���8��N�ί��+�9��<ۣu^2�#]���{G[��!�: 4%B}靍�G��z^��d�>p�����@�3�\p�7s�v���xz������ͦCzC�����=�XZϴ/"|[�dF�v,�t���عF_�_��L��n�if��5�2ު��C6����s�ħgQm�nm��)$�e�t��g��A���у���^�$Q�"��;C�ۍ�{M-�w��_�=��4�,ul {�8r��5�?
���{Ԓ��͍�;?C8"�>Ÿ����R��꿯K,}�<4!SDV�`�#�:4vIc%�O�
Q,s;&d雭��SL�Xi�ö���8vF�6g�=���I@��l+���/���T����4�'��.�� \�	If	�|6ç�Ȏ�F����XG�`���/�Z15�0{�:��UX�[�e?r�JewZ���@���3�_��2<�n�S{��m6�Af�	E����ߥ�^�C;c|tRT/鴟�q>���P�q��t�Z��z�XL��c�غe�vɣ�RZc�f᜛�)d2�p�Q׏� W�B���5K|��#�L���F*������|kKj��N!���n�&=�`��X��oF��v,,�����mN�/�Q��dH&����B����=|T�.)�9Bf���S�0U]	(H!�v73�E�߭9�G�_k�Z���X�0lU��
�L��}�K����6_���E���6�~D�c�ye�tf���p�P���+n��Wj
߶�к'ac��qλPC��� �?��,�S�X ��Ai'��C>Vu�8�K��z/�%��8𵫅�nw�EW�3��f�9�IP�$���Go�/�m{o�����F}�g0�)�k�c�åLEP��GW4�;ry�D+S�
��7e��8_��b�Ry����4{�_k_��{�B
����z���J�l0�]���-|/��x~?A�;�^��~�(	�F�z���G62�rͦ��;��g̭���VN��/��h�o&�d�^��.rz�eo���g٤sM�C�2ή+Y��[J���t(��=�)y���*w�PݮIMQ������j�������
Z����$�dLL|�[��*0�I��C�/��Yܚx_R��kv���}��h�A['�F������0���h������Z+���������4�޹�P��t�:d�:d)׭�r�c����{r��X�E`���85�gdI�����W�p�p|��ʹx����@*���,R��;jb��ZdL��Y��޴C��a�;�B��
�I�	�TO���>��ߩ���bY���mZ=��	~�PdˇX���4s�ڼ�w��{��X��f1���һ9o�3��K�岨U�
��T�� w��Qv�dg�.'59w������������:n��y�jA|<�fg�)o��W�ʙ�.7�*�j�.j*&|d�w���Yb�R��tF�s�o��Ů[3"��Cv�_}����3�X	a}�C�]��� Ï�+��(�|�����{#i��]����g�.7��i��^i�	�@Jiwf��O����n&n��L�]��hn�
�z�`��#>����k�ciI�	:��-��9�(|3}'�����W`�~m��_����� �� DS�5ڣ�;�ö�(뽅��׋��}�vYHv`��n�
Pu�[�Yr
�g%FF�T�{O�����@�+�������R7ǁ(���_�C3p��>T��t�P۞�إ��Gc.�I����l,��a�z�"��A�R�Oضv�|{��B&J`���O��K��KN�������8�� �t�q���\���U��K�Y�AF�?�js[=��-}���Ne.T�?�q�i7��xEZv*͒7	�'A29�c�:m�#�#�)�vlշ����ii�&c���"��M2��@� i�,�3�T˯���*3^�wJ�ė�[XT����'G�M��C_��wk����%u�{_�mP�r-i�!`l�k�|�s� �HK�  H�o����������u��w-�ӬE�3ya׆�z��^&��,��U���6�©�"�m�/�Z���L�nSE&���~�ʏ�g/0���)�-0�s����Uʶ�އ��aTf�ȋ�9 ��J�A�ݸ�%d�Rt��S�"n.M�a_�R��B�i��(�GG�~����n.�Y���YmZB0�@�����О7�a2�Oȕ�ّ̅��Q$�+���%�8�6a��|\�X��^��K�hՌ�s����8dI�F�>�DmW�d����^7o�41.1nf�v�TJZ���>��Mf�H�I�Y�@�|2N7Zp�I� 
_�>�2�a�d}�!_/�B��:]�<��վ�W2B��.I�{�
���9X~��j��AWF}c���uw��p��1�Db���9���eb9}a�6���l�<�j'!'#W� �l�U'��A?Ԇ�>L���P�|k�~��b/&���I���g�lZ�-��yw�:���`�T������{a���K��g�'���o�uMCa��\��i��C 
����x�J����a��wȍ��i���.�;��	בi?��
������_qњF��m���^�\Np��ثu����D߷}�-22�K��	�*���'����ђ�4XVw/Ŝ"r�[����Y�tu+�W��|��o%���ӱS���j��(��X�Eu��1!���m�W��Af�f7��,���&�[oz�W��L�o��g���+ߠH�R��/����䅰o_�s�����0�q�V1-����s竿��z�p �[�3D퐥G!���k�P�v��n>k�����1Q�.��QCԖ�a�Z�#��~U�R)���Iz�F'=�/{C-)����}'���:�m�؂d�f���&
A�l�G�u��i�M��U"8^�y��N����Md%C�g �G�
��E�V����*�Dt�H(��ɞP	�l�Z��K�4��x	]92����))H�3�W��*g竽�=�dO�������V�,�م��3z�;��$8"y��_v�v��%��cv �gsr`���/�sk�"����E�����i��Wv�A��Ӟ<_�#��_D�mӵ�oǣZs$9�9�qcW��OZy���~wiae���D�4��MLҍ��Ѧf����3b�&�oj�^j��kt}U�ؖ�3�ݦ�Q˷�)��P�NN�g\�����oTE3��%��d3M������tᙓq���|�����gY��%�Q���N�����q���j,�H���us���,�	�4����k���3
T�p�����/@�)�i�V��4L����0�ȱ���4��ɹ�7Ebvsz��J^R���/���IHp&Sy��"�f�Uj,�T$_��1�P���X*����#dBl�	�]ʬ�אez�3���_��(I!��YT9�
� 	�V������ ,0籖I�q�\0QF�E���H�q(e�u���9�8��_I�N����H����SE6m#����?{߳W7{e*��V��tk��R6���<�ow!<�,�8��L���[6�Z⇆�OH� c�n�L��[�CZ�w�Y�Z�2�%T9?�h�෬�3�od�������Q��T�^�p��:���������t0 `�j�fCtA�x��Ĳ27�f�%ɠ�n$�c�����;��0� �@qo�#~]��0��
�G9r���:���	�;��~�b
'Y{r)	=ӫ1Ş�]����k���X���^kw��� kn���$�$������k&�2K��.��	�@�U�=2h&
��Tϕ�nf�u��Rc%;�^[��Hz����F�����VWKi�%�y@�DrH�?��LP�4u2k�^��������a�r�\�����~�K�dF��)�%���e�떯f���tZOi��U�>�
�Ua��\暈�Q��@�ݧ��L�ZE���yaSн[CS��]2���a�O�B�e`7=���=Ɣ}ՙ��".� �v�U�KF�ս�W���&R��,���%_�U��6:���'e\��*l��]�7�����@m��7{S�k��c�y�o.�N��/4a��&@�4뷃�9��Ӻ�V؏V��K�{���5qY|Ҕ8{�Z]+3Lr�7L�"3���������-Kꗖ �/sa":ÈA�՞�(�8�xگ�oD�$���z#v{{Sba��:P�a�@p��#�v̆�E�l��y��6h�-�oQ�08*N?���d픉�b�"!����3\Mɫ1R����x��D��8�q���w����o����k�/�Ю�55��֧RϾ��`�������Iʖ�lHgf��}�5ϝcs
��ۣd#�
%A��hisgj��󫘔�ڳ��ƒK���ʓ��@f�nm43��\X��γ�w�Q@�j^|�+�u��5$&;�!�1/�b[���y�]bE��~���w�O5
�D9B�i�����f 1����/KJZ���w.,�(�	?��J�����Jb!yv'���;Å�(���Ψqѻ&�>�W��ʍ��YEEl�2��i��;O��S$���gR����b/�~6�S>�}&|o�%���� �_%a\I6�N��&I����O�U��A%�w��f�W�, �wˀk�g�jy:����ԯ�	�A�`�,���Q����>%lhp�5�����~�<1�����G�B�+��r8f�.]��!�B�q���!�,���E�j?m�h���q��!T7�?jd�ճe@��;9Pe����pw/���/�b]��TLO߿Q������K�&���X�rfJ���)a�읍?/����"��,+��T��J��)��+�WH �C(���n��gpN�C��+2R+�(��M<|;��@:ئ�������y�m �zF�%�Ff ��Ϲl��h:��ì��@���_�mޏ����)��߼&�z�O����rHt�k��u3�N��V�-6�� e���ʤY]�cxJm1l]b��j���;4��UNiB��;�n���c��"�WM���f���͇Z�_��w�B5�'Y~лZ���I֓��'�O�@K���:+�&ltr}�r���%�H��Q������,���g�ł����t-$P��IP��mڐ�0���<XTΎ�>l�q��8��g^���\\<k	Z7�����R>6��hWN⊶?�p�9i�䷚Ge)�K~����4I�z��7�ow��5�k�H��Q�2U�	���-�v����"��%�����Р�tK���l�Q2≮~�F:�-4�
�$`�V�*�?ܸ��%W,���D����
�i3���i���{z�vıO,`���s��.G
��`�6�����⥫X_y�����Ԑ���d�*���}AOV�t�����4l�?J�h,�Y�č��1yk�'��q"I�ii�(�`"Q���$�R��覆��:��t�vO-��ysi2:�������+����@�fӛ^�������!�mH����/���?��x�,��ͣYg�\JV��B�D�ۃ�8d0Ŏ��@4��(K3ס�ixC�u ����o�E�l��e�h������	��)��ވ|xP��='J%�3�����k�!��K=�W�_6S�`��\��� �՗�?h4t�yk�s�.6���7�r��ހ��;ǎgN�K  @��$�z.��d%=��ҏjҸ�&�&o%y����]@0S@���)Uj�voE?d�y�;Iy;�pH[u�?��� � i����:�t�z� cW�y������Z�3���S���/���t.����.�J��t�G��*�j���Y����/�G�>-�%���1]w��]Vi	����7�p��ap�ŗ��:��x�w��ԓ9�����E��v�R��,���d:ҁ�$���O��K���5)�����?���.���Լ���@c��';.�E�;��r������P`�q"��L6��z��&��k�L�g,�ɮ��]X��u���U���b��7�݉7p�P�1�;����5��WBؾ�(���w;��}�z��Z�u=���M�eHw]�݄��[��З�κ��!k�C���y`=�P��	[�x��16mIq]���ž]D@ u_D�_j,���i�m�X�(�b�]�>���5��j��e�;t���(mj7Gy`�@�ӝ�j�۹Y{����'�����)�����''��R� �3Z*(�0���q��>
����>��9�i��!���Է�}�*���"� �I־�=��Iߏ��;��P��;��Э�.�W�!��ީx��ɮ>}�4�3X�i�~%G�a:blU��:L���|]d��9�:���d�aI�<u�\�-�����X��V*���/�o_V�a����O�Z���y���[
*��B��P>T&��߄�K�#8�f�Ї�+b���������x�����8 s�4{�c���ӱ�L�,���Z�v-�6���
i.2d���!�_��i���oG�g���>a�'�
5���� ��s0KY��K�j�����DJ�*`�^(h�4<�L�;)��h-�;���^�Iß�u�>���|�>�J,�rc�~X؍���k��x�s���m���VA�7�0��kHz�ka�<�sNm�R���C)���r���HMK�V=�
1�;��܏���#���/\_1�>&DQ��a
��]��UK�1���%�e'T�/�����k�P�Vye���MXc:?�I2���{��N�f��A?�/��'�a܉��*��&�ۋ��᥇ӌ����)&Yk�`47�G�I��X�/���dT����˵���XC��O] �ҁ������n^V3�'��)/xX�=�~ �R��ppA^ + CP+o$��C�]_u�\��^��|���%���v�~��M-6h�ɞ�詒\�ŵE)Ƭ�p�F[��F�mR;�y���K��[��E\4���F�KN�����f���ا�]~�3�Pކ_�>�PvsP�Q�I�7�H�����%���'��w�~0,�,�Q�m}�T��+J���r��B��!K�C�?߫ 3 ���bi3�gL�K�~S���c�| a޻��g`C�U��q?(�m��F�<nX�&���V%�R:��Q����� ��ݥl�S[;�k �2$�n���E�L���[�I-\|P�7�h�( S�~��~,��냄1��8~Ӌ����( �4U�R��0��EM t�|h�@������*���g��Q�1l]�e�Գz�N@FK�J83b�܍��h��x<�i�v��kW�lv�t�ܨ
m�m���{��,��E7�s��]�v�x�����]���2F���m.��#��Ғ˹����ߡ��T����U�h���V��Z=��O��yڅFiW�C�56W�>�ÿA'AI_���x�B:D���.�����l�o�dk��ꗚ�%�Ʀ
#�$H��mQ?$�	�������1�0.�R����>S���C���5�a����O#%U���i%B�Ͼ��k�ş�W_�	���K=�o�V,{?A���@����d扃��#���k��5��|F��{�=g� �0,���t�e�IB�d��G��v
��l��`�ۜO��sX����D�K3��6�~��h󩭈�����Gj��W��p,�S���1#R���
)z�d1�֠��L�M�R��2�_�\�����aj�\)S�~�o�� ��D����ڴ8$O�	6�'�8����Ɂ9 wtߝC��p@ߚ�545���������E�C4����uw�.�b���!�酪a3���Q���d�\��qt�_�J��@�9���>Bu֩"�ǖ��%DZ?�I���������)Ϛg.���.Ų\��
*�x��xwE��wt�ͅ5�O ��Q5C@��U{��%���ڸ��7��KT}��v��!�`���@6��58���3����j�T�/	;��v��4~��˲]w6������Os� �;�xT�/鏒6��6�g��N�-��9#�NŜ�]c��L��
O)�N��E�Zx�E�B6���A��Ĕ�U�)�{s�p��\1GJh�5�c+�@�
��w?�����v�z����="�� �5H� 	k����&��j�]��Z����T0�O��x8�6��������we���D}�j���f�ZӀ��O|�K.k�nc��X�mU>HOKJ�.����6�tN{�Tv��q=� C5pW���#}.�c5 �p&�k[$�c	1�w��z^$�r��P^�, �ͻׅT��O���]t/ J{�T�*2�÷�V���x�<��ޕB�3�.Di�����u��w�X���F]:�&��Dp����h��Ȧ}1ߪt�M�H�a�Q��/ܶ+�ё��N��-@pt�V���o+�����.z�1pa���CW��,�}��o��p���׍(ƏF��~�ŋT�z@]��Un��.�,z�-.�AF�Rך�;kT��5�d2�"�O [�xn"B�_�$2�zS|����Vp��,�$�k�g��/�a>i	:�ua��5E��"�ๆ4� �J��^�:���u��;g'}�+�V`�G�����|�ׇ��[�n���]��x�!%Y~�J$ӆ��v{��`�h�lyRU�(��߮�%{�úf�X?�0ٚ�7 vѣj��'��YT��B݇{�?5������+PP�*����*�Gj�_0�MPO�n�K+�ܿ?� �u9�GN8a�d���N�����S��S�������L��D{�ޅ�x2�=+�ae��B��|��:�u�=h�)/�ڟ"ώ��V����Q�$�]
��F�G�cՒ��`�"B��|��Շ�Kܜ�}%̞�G}?�T����,^�f�yʺ�KXȍ��7bW�߾iװ����Q��`��|��Nw4H��6��m�.������H��ou[PkxC]d�Y�5@`�Is���PF��A8�yO����x#����e1���q����w_srU��W($�<�JՊ�
�+�y�T��ajS~2{oV���TZ�d�_&���|EU�����T�f����U@����z���V�/�n$9�)S�J���f�c��kz�5�#]�Gȉ/;���9p����h�&�1��v�ik6��C��T����.B��E�,�;s!�1�-��6R��n�]
��w�[�N���5�ӕ�%�g�X���8?�ufv	�����_@L僡�6?j=�� w���Ir���\r��9����GJ�����m�~ׯa&���c�W19g7�}w�Vc~L�~��nA2Exܧ�7�-�5nR&A6r��2[w��w�}�S��z�yՆy\tȟ���SxG�H���=��/b����91����Q�f5��<Ey��Ne%%'&�Hݎa%>�J+�raQ~� I��JʪB���(�����x�[ŕiTUU��lc��>$����;6[�����d�2�'�'�y+�=��jzjjUm����ЯG�R:�'ܾ(��gzg��3B1�f�h)q���7��˥��Cђ2-J<�Xn��e�Sb��'V-����in{���*���j��%!Zn.������5�O��0�;�U���x�T�4`@~i'�\�E�����iJ�<�z�ڎg/[L��.<��t3�U#_��ѿ���&��;zx���e�u}~T�p�9��Hʨ�����a�C�d��%��_�'�+<
�8
���cMRj�]G��m�y)mٴ�_�ߪͨ��;���K�>��b�UȤNl�i�<`�k������X���l�Y��ҹ��`3;['�`{;���uP�L��?�9=��Q`��jH�+F��D�^M�v�yq)T'ey��[�L���u����3x�(.%���՘�����V�y/��_�^�����;m�*�{*��p�ø�yǣ ����n�4j��)O2Ne� l��9^����>'�w3V�5G?E�Vm�5l����Uv�,z�
y�r�M{O�i�h��{�����9����1{��R��6a�Ռ*���'�o�4i�$��^�v�V_'}&[�P�[�ã?+���$Ûؘ�L';�]���&I\S�%m�����b��y�	=u��Y;@;f%�!��;M�B�Vs�v����V��xV��O��;]���׿.�����g��;t�p +�'8�C�k�(o�!�)З;�z���[-�X�6Ɖ��i�rsaQ�-Q�����aˣ��_�ݸ+��˦U'+Ob��N���)t���<�ƙ x���,�4+l�]}k!\�Q}�Dq0�궧�K�P�Z�΍�1��xc�iS��v��+����xX9 -}.�j����?�� � �o�{]Z��5~��$��x`@��W��N�?��2W�%��GSF���NT0eN��w���TxݭXQܗ�S���Q�@�4V3�2�+��+�j)����W�t��h���4��8��AfE�Sވ}&X��Tbc
{{�$̽?��C�:����x����@G����2Sށ�U�Xi)}�$�����CQ7�K��-f�M[�UC��A׊J�C�S�S�m�0H���������ߟ��E�����%;Į� ��®��yuǪsjq%53a�#���&���. >�[����;�k&~�<~��8�����<��nY��n&�׉�'���N��q#�R�.杋������B�ki MY� N�V ��0fJ����6��[W{�S}}�W�X?��Y�k��z*#�< %9N��
ѯJ�CUa}�@v1s?�P�hU���� >*���ě���&^�U��~�3��r֥�ԙ��� �B/1�?j>����_.eK.���V� ���>�O�"���Ñ�U�R#��Xnϴ+zU6N�)�m��ɖ���� �N�~�;�Bd�{y٪*�+mL�է�|uB¤(�-��Y~�֞�&���g� ��Z��y���;�\�|M�����&����ԥ,�4}���q .�[�RK�:@��y@2��Z	���,]�Z������_~dj݅d�8��jߡ|��4���o�xA���C��U�-Ȯy6\@Q��R���|��aӖ��B�kݲ@3^����J��x�~d_�>�k\-^�U�^�J��o�|9U��$��w���ɔ�����[
w���}� �T;�GfM$���07M���~�E�k�B�'�]��\^��3�ϰ�uOƏ7�V/7uqܙ�ö;�[%�, ���ʟ���(�u�%m�;N�L|x!V�5��)������ֲ���u���M
�yI$�0�_u=Vm���_seک������r��`ՆU������m��i�n���tcy]��{7��l�����7���|r��QNN�؄�4\�xCM��g?V�}��1��a�O�m�;�n�iz^�u4�q�Tyh��e�t�"�=���0 �#�ڀ��N�P��+a��vG�\�~�%L�u�&�[�EF2��o��~;��)���.2����+���<�q�}�I�i�bK�L��5к7Q��%<�z��A*����4��4U��|��a��9k�NӬ�.��H�X"ŉE�(�����PZΡ� �'!�ko1/5j1�ک��YP��<��D4vyc�H��1]���bk���]cO7���;�zpПg9�M��Wo԰E8��H�e�'$D��W�����K�z)���G���j�iI��G��^b���������1w���@��;�y.C�O0�v�;���h�n�Qk�a`fs�꯭��Db/�W�"�M�?������议=�	�1�z��a�s�g�L�'7Г��G#��s��aI@��`'���/��]�]���vfƝ���1x ��P���<͵�3�B\]��u����6���s�	�rb��ۤ�������U��'#����X���s�)���>��y������ۮ��V����h \4Z��E�&	��[�Z��K����#��c̟ޞ�w����J�_O�fF�h��j�c���7w��"��]x<��jҜ��'Y5M0 �sMO%	������e����kT�AUx��o����}�$�b���N�`��co��xD���?�	��_�|j������7ޣԐ�M����b�@�?��%r�j�M����hbZ'{�\��d���O����F�OG�y���8y)�O�5?�g��z�0L3����iݹ���˝`C婙��j��_�ɫ��ټ����{��n�`=���:�����{�ࡖ�jJ��ˁͿ�v��캆�h�6��]AlU��V�Sߖv_������� �p`T���M���|-�w1кa�dd3�f����/q��7��Pe��)8
�I��OG=�Y0RQ��P���Х$��U�4sF"�.��=z��;�̈́����ۅ�30�c��?ܽݜ�5y�ձ��C���#U���	�����qm�ډb�Q{�Ȝ���w�v����RAyb#�>�6Mh���6C8|t8p-�0�d/G̞�Ɵ\�$X���h���>�~[���
�]��&،y���GU�xFT@Q
�d���p�A6	��)���_�a3ح@�;��1�>*�j��M�Q\�t$�G	ss���n��Qu{��#��?c��^3�;�Ȳ4Ҝ�,ڣMʕ�V�ݩ�����פ����nnD��o|��)<{Q%��{��e�i�i1V��c�����䕮�U��z3��]��S�ƢA��J��S��@���m�s�B�Q�f1&����J�1���Lv�֓=}ڥ5L��3�u��Wi�hR��;ZԬ_���0b]M|�����n�_�����j���D�H?�^�Q�N�m`�^^%%�����?��9/�@�5��n��5��f��Пaj���g��,��w����ש x�[����klщ4�5WdQ�E���;��( ����l1m�=��/���wf��(���x�@�o�� 1�o��NQ����G_�˭��&�8�YVp1(x�KO��.��]���	�m�S����ӿs���y~L1"�<~�~Kc�#��b��W�DH��z��$�#���ּ�cn�V��:���!�g� �:8v����Ӕ?�I-�$+ v��s%߸Π��h�KPL�#l��{�gos�[ױ��!�U�ӈ�G���)]����N �Cu �I��������nB~q���%`'������e�bq�,�&��桮��j�'A^i`���h�ub�%�.�'?!�Pg��#�I��/yacżJ'/nq��/s�
�I<�B�ȝ��[y�?/"�o�;�s%�23�O6�粒�'oH��q" ��EA�������<�����;�`j�_};p��|��a_L��)|�� ;�u���taM�mU�I$�s[��D,�03aKt���f
*B�kE���?����+���b^�/����*4I�HHšH���pSE���#�����ͅ��m�����j ~�ݎv�rEt�#���x�W�p���ߓ�!d����3-�0ET�Sj���_]�4�|`(teL�hu���4q+���K��̎����3��_���w>e|	lX1r�=];v�A���zo����b[O��?s���K#�ڞ,���`,o��}Q�H%S4Bq\�eS��	Y:�jGL$��D�c�"�x'H�ua�4�_Uk��cmg �.�a�Ɋ6��8��T
B��}�]�	�Q��	T��\�PͲ�'�"�B�f�KX	<:&��㦍9�a�9�]M����m��y��+���Ҵ0��<Y��T�M�0�K���Y��Aj�4kg��;M��7�+Y-�Y5x�>'��5�����B��P_�������b�^ƽsVM��TSn<N:@@�<�U���,̲Z,��n�{t�k��P>`�9Pq�|>'/r�W$Ϲ�F5 PԸ�C��8�Я��nF-�CrW1]UYM�q�jG���gGT�"iD�w-B� K-���gW׆�D�hE8B�̗��N�9K6�jWۀ씚�����\q��RWخ�jyD�2��O?����m�n��E�@U)<�:|w���JH�HϢ�@�X(@Pf�v4�vy�u��j�����:���W�W��+v|�3jE��>�5fPh�M�1�?_��o���9
>�;�+N���?�;��ݣ�'&����������V�4�ʓǿ�ϭ�0�m�s��>	�}/ H���G�c����[�:i��ve'/бOax�f&8��Hd�L�u�-9�qP���e���Y��2T�!9=�z����R�x�(>D_��H	̫~Q(�W�4�?k�V��Q;$0���#����v~$�X�~�u"u� �6�O�PRӥ!�2`��Zpx��T[�� ���+����a@��K��c��DL*^�]]�Z�m��!M�g9�2<S��LO3��j������_�b�hO˟Յ�J�����ޖ9��@^�T�@&��uD+���O������ �ۑcX���@����`�,�)����b�@�ؓ5hgM ���xX\���7#ʓ�K��3g@��q��)j����|�RJ�!c6�c	ةuL�ο�J1�{��؋A�Ӽ�ߋ�eIuR	�I����gT"H3#�=�!;���� G��*����_�_�/�d�����?o�5��j��J~�9�j�./��2�9���&bA�X��z"���.�{h�ۅR]r9{�_i"���}�J�۰#�����#Ӈ��	��Z�����)����+.!Ƴ8h'hw��VE �)DD��~�Q������&d���@}c44���y�!B2���Xr���Tp��z����!K�DKef�w����:.��k���*"!R
J����H�R��0���(5�*�"�1����H3��59������������Z׺ֵ��g�1��j�`g�4��$��*d_�v�+�M���S�_���&���,)���\��������5�C�Jw���v��כ�yT�U�`��{�&h�a9oP��v8<��_Y�O���@+�wӤ������숕0o��iX�he��f��M�?^�$x�"��	S�An������?��3/ѐ���G�0HȨ�
=�'�̛. ۬N#�n�j�¹�AH��q\���!th'_ǃ�K�OE�g�Q* �j���:��t�^`��]a�+�m���MD�A��l�q4V���}����������j���+��7�����46D�hA٦���U����*W耤���.���[{^�BG�Ô�$�>�1WU�Y<C�h#꣤�S��uf�4��Ƀ��6p�����2����hd�yf} �6�hy�YHR�ۏ��s4�
mH�n֤RP���6�[��,/���D�y�S�{�2�}�����2�Ě�e��D&�ȅ6rīn�yKb]N�D�D\֚�60G�cYn	&k��)�	p�ι���l��ڿZY�,�`�`jBa��חn��WR߁����&T��H�!6���@��4��]s��\��S�)4{!hS���v˾�"�����GBS�A��-��W��?%��1B�02�`Y��{v�/�5SQo~�����_Ǌ;�5�@2�G������W���ͬ�='��P	M�_uo`�W��u��4�S~�*Z'L�OMR��_:�\��3]Gl���r��O��ǌp�l�E�k�A��*���>�*��Y���\F}�t=PgC�~V�++0ph}B�o�ľ��y��?��*����3�G9���[*a�\t.ߦk��0w��@QE�}��3������a}��h%��o-#v� �e(�%���D~���M�n9�A���DO?Jt�tV��wl����O���f>���j�u�Q[�`o��	�J\[��C�?�y�ݠ�w���"�L_xS;Y��B^<h�g�s�E�)t%����Т�Y���d����W^��+��=�$� g�uɮz�鵻�go��y�Ys�&|V�\B'sx��܏MR����j�䩩'�g��K?kTR��g�7ʆ����1�?���݀�Z]�ow fzM�jwt�XfaYz/!3��̪7�z�H4��/	D��g�ӛ�#5^yʭ������}2���������,���Z'�$ѡ����Jy8S���6V�7Kr���_�_q��a8�o[T���Y�vz��ThA��o�8�B��wQV}��R���M9�s�<+6�d���ݗ����8)��[�fc���|���~s_
?�q�Nw~�T˘�&R5�F{707���m���֕lPzk�[r�N���F�C�`���6�Cޥ�S�-1O��2��B;���*ɩ�8�@x�6����@h�I��F}YL�	���{�����M֞q���ER�&/�]���Guƻ�c��U��9V"R�x�ӡ9e���-RX��=�4�lmU��G��K��T�35�8^7�q[����dO���M|�J����P/*�9Ս���v��"��y�&�f_��f<;ɉ��>��c�|j��b�<ٳ�Z��@ؾ�aW` j�t�|w��
��B��+�#��L����jsq�\ZL;_��hf�^���'�����Sh�ȱ�!lB4�������%�_�w_k[0P�A��7�L��3/;h͙M�4�p�����+�^_�����j:����]�o�Xo��e��d���z���Y��x�
��AYl��=���4�VE��7�0�-��^��Y�GUH�9Y�&��ճۨ��p"q'���M&=L�>31��!y`p��0b"�aH@W��,me}��[y��HZ:�=�C�j�;�����n��<Ͽo��:Iئ;I\Y}V-��>-Y�F�'o�{�Z@�P��1ʝ��Z�{�ٔ��>R<�]4=���@�`q�$� ������][�.��r��|��Ķ�����UDAQ�͑d�9�<M22��9�x�|�.��������~Bs���;�+4���P���
�Ƽo�i�!���{]i��V��Q��
l26�_��$�kw�9v%���ڇ�C�����TTt�ӻ)4�$��S���oWΩ�� 7��qgv�ͩӔ�)�@+S�[+ۭ��k2|�0�kӷ0M���)%�s�gM<~��n���32��/��nQ�_<z�!�5]��o�G�ƴ���%:�n�������3���=��w���#��l_4R��X�	'9�&�3,��4X�.q��cN�����R����X��О����\��h2tgܠ�i׫̈́��v��)3��8�"�z͸�{�y��'�<i	ƭU
�V�*Vj9yq��}I���	���lL��n\�S�k��0^�
���i��xP���%���@We�h�����j����Q|�x>$�N���Z�w')�
L���G����\�
�Oٙ�!|�3��`�u�X\{�h������m�� ER��kz?���~�R[��2��N|f�頄x�`�����B�ϜAn4\ʠH�t�`RЂz�"M
q����N�s?�S���}����<�dq��`��(?{����?��{+ʻ�����ؔ��ZB�7���]͞�j��~!�����w���h���w��dK�Y� *4�z�U�جT�%�Z���_���
�A����`��s�o��q����,w��W��4�9f%�Ŷ��DPx+ͨ�:�r!��#�v3������,��Y⢈Ec-TH��^���	��I<��'�gz�t��h��p���͍����;�׭��&Wʦ�3,��j��w�JTr�<���˞�!���iMm���R�����ߖ]�ﶍ~z�E����nx9�����)�S�Cr��>��ǜ�Z9���s�ZfS	N���S�P��a�zjm|*�װ^dv���9��x�9�9��/x�U�	"�ľ�&��K���&��y�T�	Gڮ��b���~��u��Y*)�ܨ�w�����K���S%ߎ^2�gsG�� ���v�Sle;ت6��M~VhY��Pr!F�ˮA�/�3h�W��hiT��I��o��$�]:�CH�v�����91~Y�K���#ô�X�_dCz�-����#�M���R�r�ގ�W{�j�9�&5����;���jR7$�#�ʞ�.|�I�j^�������ņȔ�l��mE�Mo��G}������Y�쾠��1~�
�F��O4�JyJ��[1�CĠ%�fq1�u�R-E6?{L���6TaQ¤��^�T����@B�;p�o�5��ߍ&|��{qw=�a�W��;ǔ��26J�!U�Cb�Wk҃�W�j�� G��?:�3}�Y��nJ6�yQ�BU�?F��J��Ƣ�w`�OQ��Sz)�2vfojj����}	 	fi�b�C�9�e�]t����՝��PNְ���{<��h��?���|��|}���{(���� fJz��M{k��h�[�p��i��H�r�X�Mܒ�_ ��)4>��P�S�)k+f�0Z^�)Xܼ!1�\)���|���6}Wԣ%���BQ��G^m���� ��Ge	�t�wb���/{��SԤ�%w+�/7Ɇ603Ngi�z	������//�m�����uW��.�=ϐa�����t�����b�Cb^�;��K�.�Y�ֺ��ɬ?M��"%���~7��a���c�G�s�^�G�ݝ�n������i�a������6O�]R@���Ϣ��U�i?��������[h��e{��x�c�0�+�S?���'� /���06*mą͜ـ[�! ��n��'BxFV�����fxQ�W��{
��Nxf:�����g �;�\�����[��.FӪ�RW���v�'}ʕ
�
w��;j��#%��y2Vm��	��)��lN��?g���r�u�e\����R#����ڇ�c��2��N�>r`bb��G�����0%\�]Q.��u��G[��O��v��/���k��N�ܺI<�]%�	�_���jV�霪 ~>'e��fdX{C�K�ӺjD����yx�ޤV���
���,��ܺo�����t�y���V�d�����Jy	�	!p��Z��/��^6����R�V�����2���u��qq�"���?�}[�ﯲ{�.�ȱ3i�P�g7�ؤ�� ��c�h�:Y����ˏ|�kht�;�h�UeL�#4�V�vwOd"S%/�U|{@�<^�՟]O\���M�҆=�s�Y�_��30O�J�ϩT.�վe��i�dn�
��T6���j��K��M>��yK�Ն��l|Qf�Z�j?Ea�)�=е���kR�@wS4A�v֙��0����� ��?���2�����C�m�&t��o9���N�A"	�ϼ�^��l;	ʽ�M�k�c�rU��|���$��&|̵�c@ՅI�\h�;#=��N�qU6��~�e���|;B���|�Eo-a��w=�
��
I�"�T=�X|�����D//�~í���}I����R�Q�M�g��w�mA�/�����-��4������؞�ӽ�:͞CR~��e�[ʠ*͑a��EH
r&�t����3��ө����0���o��
>��ŕA'��T�jO���>�η�]���U��m<�_ZEB���n�Kܴ�"�� �aﴫ&�jJ��މ�v�l���ݙ��x�Y�+�6s!��>7�k���^��}E������+������[-�t4��tQ~G�GuQ5b@���Y�����;UƮ�ɹJ�y�����Ի�Ei�Ѹ��v�#�3��z�ȧ���0$k\CIܒ���1*�W�hדF�g�hrq�N	� /��:��`5�=�CT���!��Q�I��X�O�LSY�����Zhtr�'(���I��9�g�T�:|.�(}.�tJ��N��祖�g*⩟,~��gMn���i*��a��~8j�u��t膁���%�;�ZQ���>���s�>��TY�ʼ�v-6M�M�5��t{;��=�ؽ���>��aH��$GiZ�TV�C���KC^��y�2H��ܯW�"H�3�gQ[�!��/9��TL�|X1��H�=���9}�8\�ޒ�,Rya�����b4n.�	�CŃs�;����>s�-�@�^���2��v��YN�.�{d�|��m
+l7m��{�ᘍ&�j���Ǌ�;)q1<���;wA,*Q�%������bȻ'I/��^���w�L�@� 9�6Q%�͔����Џ�Nw߿3��\���]������}�w��K�!�>Γf:o`N���'D15I���,t���-)`6i��B'���ǳ>���?w�ն+lW򄮫�&�1���Q�	�3�p���;9S�m��M����mր�'SAE�<*:���$%� ���8����m_[��(˟�>û;q�	{�d��%&�����O0�#�Dpۋd%e�YR��S�Qd�}�8ja�qLm�|���L��Q3L2k+�\Ko����R�=�U�c�A�e����lġow~TT�E�㾘Fx]3�_nVd��PHx���V����'U���$�4E���0����]Q�A!�5}\L^�n�@��������a}�ϨN�p�}����	]� +J�\}����m*�����d�L:�:�)/Q�12��|�s�'���g�s�7��E��c�=���Ϛ��W�}�?-9%���:��T#;��h�zz�_�:K���h"���^�}�7\�5Fn{�x_���J�(e:+�-R�I��e>�a�)5\QU�M��v\��>�[*Ԫ�^ d��T�W�^H�(@~��|+���oe����}�ͱ��xa�؞����c��X4H�*6��T�<�� =Kw�^����|jE1�����gO�@!���_jK�kLD!�jw�Yc�MloM�W��m����s��^x��;�P#�μ^����N��aO��r~���w�K_�8
djB��Sk-�<�=,��~�K��&�vfc��5��U�:�
w�61�5��y'������`������QUO�C�al�/�m&t�G���x�J�+|���`I&eo�Ͻc��H<��ʷ:�H?L�j�NVx%I�|	�jJ�ZK������f�̢t���r��4��64P0ˑ�9l^xq�Lo��\c�HNPn<k�����{����Ť�f"��],q_b:�M��)�
|����a��aVW���qe�]��<�-�S����%���������j�g�
?p��S�ފ��B�+e�7J�?���<_JF�u�c�6Ka��=��$��S��~�.n@Wp%��gNN���*3r��|�Zȵ�1��=���nvK��K�AYbd�A18x��K]��Ix��if�B�p,���w3K� �h��<��3�Rd��A~��Kt�3C�B%x(��X���`�^M|}<+ ���J�(�Zlw��)ͩ�M#��}���y_�P0�9?4�=g��"Ӝ�t�����Q�f�N�l�����ė+K`o4��EW�{�����H�� W��Gd	k��?�CO!���1��zt��ϼ�$�D�����ѡ8����n���Y#S%I��+�+��ysI�JҖ���U�3�;r�
���B{�}X��2%����b䝣Y0�,�M�aLP*�C)��-[$q���[揎��9�]X8G�Ն�w��,��e�k+��ڢ&$Pռ6ۧ{�~C6�>,8�^�_Ϟ���b� �W�)���j��~,t��q���B|��S�V��ҫ��FY}\9A)���'��g���^k�v2My)����`�&�����2A��7�9�*k0)">�&��KY�>�v�n3�'v�<$<����dw1{3�\��_�KQ	4�ޘ��M�ޘ+p�oJB��UJ���8��ɕ����t�JW�GC��p����<��]?E�q�c�'@�Rt�"���H�۱i�D(�N����/U��\[��y�B���֜��Ѳ��8jpb����K���>+��J�箻xlg�^�Ӈ�Q��5��R���EJ	��"�j����o�)Ooq���|LDÈ���˛}ZO��U�f�~(�E���*, 3��6[�o�����/�����a���ͫƦ26�H�}W��6���nD�M\�yt$v c%	�G�I��?Tb+Yb��=�۳Og�[�[���=���C��P�f�u)	0(�a{�G��w"t�?�	�;#�ly���X�~T?�FS0ǁ5c�ώ�Ѵ|����G�(��؛):"e�����+�P�0{�Q�ݯ{)6e	i���'�����s�c�@9�1��UIp�ݮ�+z+�)a���7��e�HӺ��N��VS3A���� ���l�9�H<�n�T(`M�kd��[�mc>J���@�nU)ģ1�D���[�����Qz��?�"�UWq�]Y.���� 6-$̌s�y ��&l�t��'�d��d���*���<�r.\ niT���ރ���{�v/E-_ۜ�|zț�³'��sz�|Zȏ�a�59�ͼ�-ȰV�mY~�������e��d���5�+4���vDTK��6��q���@d��H�wK����w�M��݅jC8h�3o9�/�_��Di��=A���r7�?�~��Q�~����\r�<�T��=*�VbQ�﯇L5���@�y��K������ ��&Q蝥�橡�-�4$�Z���T�}Lp�����;P+Ϗ�<�����{�(Q���t���ק/�k�@��=����v�1s���j!����K�_����,�+1C�g��7���?���{V4�U�����R�rS�����ɅO���Q��$��ӚR�&�ƅK��� �,���q�B�ևbA��%Nv��8"�^����#Wb��r�PL�a�JjII�2��~�y�e�̒�ow���d�0�*�2霯v_��v	�A���+A� ŌNb#,f�W�[���0�ѽ8�;G>�9g�G������,^�I��EZ�i�oYhA�rܑtI��>�7�V8���[��a�D���14�>E��Xd
���Ύ0��Y�ud�yR�6lb~]��t�H7T}��;��f��i�_�2��$1i��/YX�U����8����*��Eٙ, P$�D�˻0����{Svw�Hj3��4��P5}��"3�5��,�U����v�@���)�Em�
��ϒ��VtP����D��8�N�����ށ�~Z�*T�;m��!E�]��ȯE�I�g擟��|��ܴ�'/i@[)��F�S��̳���|�u��S�53��s]V{zgIdU�v�(C�=��*���4^�">��	�P�`�M��[?���},a��T�I*��á���-9�Ê'�\5[��c0�Z\6��!�����C�+��M����܋�`0�v�6�wst�p徥4Yr׌��J�6��m*�[N�B�;l�Ì��P�s��W� 6k�:k�5&&J��mگt�+	�E�S!���{�}�Ͼd�>[^7���������`P��#�PKO�[H~}�@�(!�>ܱ*���f�@~e)l����,�L1�ޛ����y�K!� �0t�ɨP!�fǭ<[k"+p�o�;�է�ln�7�(���xDنތ� ��V�8*�j���9p��Y����q]1 ���aY��qn���%�C�N��(8��f>Λ"��1
��=��Xyw}�G�^�WҔ�fe֓U��Jo�b�^ל�'�cy�>޽�cF[^��]ScP�Ǔ�Z�O�I�"E=�̯�~���.�רf#��k���xT�7���BRdq_N����/#���o����W���(�1m�Z��o^�~��� �Op!5�5��6r��=��$\�J݋���^=IshY�P���(�N����/���5�C@�����
�9����s3-�H-|���4�N��.­�ਪ�w�)H�/ ΃�߼�����ٛ��_��q�q�{�Wr !x�.>:���/��x<`;�TQUB�\���'�}��*��C�������!�S!'��v�cve�}��yb�[l��bK8}k`Ʒκ3�n��j�9z��Hҧ=Q�H0��7��Q�������MӣMT%*�����0w�bV^Y�I��7E��m���iz5N
�绿��[l�Nڋ�F��9�IZf��Ws`�AXkD�	9/�IG ���қ����\1n�}����x��n�1�{�O�
P٫�LF���/'g؅/(C'JRl�>M�B�<d;�(�F�����FO,wj� �>����VR�/�?�E��v�4���@�s�������Un� ˂��� ^��b����6361˿���^V���]��z�JA��t��$��7�5�fSTF��f�޸*h�����5��;�Y�1&��=�/^%��h�*���9׆N�
uޥ�H�WNj�R\�J�-����~��8���r�)n��R�Pi���ߦ)�l�6g�qm!�~_fZ��\Y�)|b�����u���%-湐�d�/� i�$�w (�a"��1�����(�VN��W�ϭ)g�Oz��!_ߟ:t�Y����K��^���#�o�P_�P'�������1m�ؑ ���g��y�����_�X���㘋p�i��ދ��ɔ]�[�Ξ���%P,�A���N�]���lL�;���	�Lb�8�	�	h3"],�g�A2��/V�肞�����#Y9%��Wnϋ���6���ʇ��U8��\10��?�)��	�����S9*�� ����Lȁs�.1�kȊA�ӎ:U�����ٶS�V����P�_(0\Y�qa�i��7H�H�F�"A���۵���@���k�3���	���]���Jl������l�9��̏�p���W]��"S�}[i���oQ&�>z�?vZ�7mmk����'�Bvk_]���.@�aa�ِM��r,���E�f���6*���β�`M�sgQ��n�}Ҝ�{�C4�˙^;���dٽ�M�RN�\;>��F�YH�4��*-G"<��EX����̴ܲ#���M)?���Wa���`V���g�O�(�c�@�,'T��mB}���[?��E�\���;�0
IC�>�����������1�I���?A◿��q,xI���F�@7�<�I�(I�n�|�w�۸�J����id�4}�J��Y���t�m��<'��`��:E̎�'���,����d���-:�����ӎVsa\j[�\���x���jg|GYyc�"�ty��|	�{��8� ��58���'��-4=]�BKVDn4Zm��=���sքɄ����<�%�h�ϐ s[MzX�m������:�XP�V,����4�]�@_����E�o$$=�rP~���qm!���+u>[��)����!5ܛ�ŷ��EVu��f'���˙�S��w���E�@�8��w���m�ڍy��|��st$ �]�f�W��'�����sK�-���k�ީ�I�������J�z��"�4xg�� �`��G<q�l��B�<�9Q~��sVQ��?dXr������w��L�'.T*�MRR�ܿo#���
�`�X��N<QD^+��?|}c݁I��K[Ǐ�7|(�L�B���#�}�T�?��R5}\�b�ô w�x��4�],XX�j�C��r^���{�W�e�q	�3��z�i�J���7��dE}v��"O����7@�����w�0���̯���J^Wi��T�b���*T��!��}st��ީ0fy�q+OLҨa���%Bs�N�~�K_�;�V]vE�u�qɛgP���}C���$���F���&���>��ܲ�@��p���c�y+QZB�����o�z ���)���Fa9d�^�Z��IQ�ñ�/���*��������E��T�`ߩ5����aeD���L�N�m}&B]�/=2���6�u�
��W��}�ʦ����T�/��|�.��+O�{���ή��U��sByA]v�k#�������XW3��+����N��܌̮�:���P!��C��5��a�����v�����N^|���&� ����*�wH�F��p���Cjg�����=�;0�CMs%ghuԑ���bcd����HL����L�œ�LB����v{�����=��G�Wu3{����$��c��1����U��_��<	��6�^��a�G���5����W�ߊqw�M9��*T�i��kǩ�y �1�W�7�,�c�t�T��;/�<x ��O4�.o\r&v�H��h�\my�5��~�[�W�L�Oܻ�)����� �|8�9�|��jvI���؛)m7S7ӥ�Z�'�IF�x������e�z�C��>�}��`�}9I%���ì�����o�g�cX3�������ؼé����Ώ�F�[��i���2�+�0$�S�fR�z���B���C�#N���zPa}�l�>��ݽyAXW���QA�_�ek����b�ˆI���+E�T�s^�/��΂�[+��������l�T�kgD�Q�N�]���=a�g��8������fP+�6w6Yo�=�#:mт��<Y��C�'��d�#OR׵�Y�{���6�oe�4I���4|t,��O���*������](�]@��EѬDPCC��J���w�ZK�F�=N8%h�x�;�����o�&l��t���(d휢{��_�*3�~�֪HUPFC[�`���g��b�7�g�<P��u�ɡv����գ�Ϭ>'$�-�x��[`��f�U�����u�ހ���Hl�!t�!k��,8`ݎ����}���W1�N(�oM�&	�|���j��\�2��iw�2�F��B��@1�۝'I���v�;N<	}-�t;.N\�^��{cA���D	��\�8�\�?�K�]Eΐ��A����e���W7)k�s`cY�ޤTR��{;�($����v�Kb�:@.jd�Pwy���$�k9e���f6s8Sa��|���t�=O ���G ���_�$�gKO
1�.^ů��Xe8iHn�|��8��]o�Ն���)��@|����ξ�><gt�L?�S@^ʔY�aT`A니n<�P��*��>�E`̱�̵�	m�2t85	��x�^Zcz ��f)
L�1���*��m���Z��9�i��!n���H4�y.��� ����'�6YD��p�G�\�X�RNI/𵪯%�Nۿ`�-���� ����:V~U���x3w�m!r[��F���eRoL�����(t�JK�m�9�M�2�@�]������	b��5I���{a�y����!��c���j��cD�@�x�����k�;�{K:2��,�"_���D�J��y��AI
E��vቮŨ"uN�`�u>�oi�F�C�~���Ӕi�&�@C��ʏ��s�T�j#��s�dK�j�n+��e��#���zo�?�=��ⅴ=x��	Gᩳ_�f(|-���|?��׮�OJ�ԛ���Wљ�$ql(�I�x��&\u�#�|�i�'jsP�y����rydXO�`���'�_���'�_�3r7�x�䶢W�K����l�5�ȁo����6:&2.���K�������V�ho���Sc=�_��Iݐ�J��Gq�������˳#!N�#,����|�O�ؠ�88�h�z?'L��`���):K��G�n�c����n��";�U�
6��=�c�o0Xlf<//%��;�}���l�ʙ鿘��å��-;��̔�2;gl��776ZD�3@7��y�Z%���)�ӓ�3��		���5_��@U}�~�r۱f��V䱪o�pedzq�2k�t85�=ԓ���T�l'��6ϳo n}������,�s�,H��_�n�̊.�8���q��7�-����Ƙ�l�wta�5ke-�P��\3�U�$�" h#P�n'��`��x��aM��{55gX{�C���N�v�UM�.�Jt&������-���#�E�x�\��\��5�B�֞�s���7���H�Ū�X$4J��B��dU8#:Mi�а�7��5Oua�^�5%���o$��3�$�$�v��� ��$m2�Ag0[a=-܄�ڝӰ�~\�+ `~��^���_4п�+�<Elq��s�@�^�3^j�k�����`'F)0�à bNAŽ���!Ry�A���=�q%xsʁN.����J����n��~�����G&&�� �F�x,	^j��5���8��Vީ�>�I���`��\��-� e��'�҂?�u��20�t���\���t%q���Q�2�,0�+��!��=P��Xn��:��Uo�����m�3��u5����3�֔�ʩ+!�������+�ak{5����sѻ6�St��mo,b�Cy_@n��vc�3tc�b���z[����t������Gb4�P����k�W�����[���Rn:���$�S�kH�*�víb7� ��g�L��𢕺�w���g?�����7��(���6�U]���Q.m��1t��
Ы\0���4�?%;Rd*21w�ܘ�u��|tC�= �pb��Q���C� �c���ێ��f(\Z�~��O*�Mn���l�3v^�C��������L�+y�21��>�:�Ƭ�<ۗ/��pW��2�� .��G�}7�l��#���/@)F<����4��}�(q���Ϻ��"h�7�57j:o"���ᖭݐ[���5��u��c���c�t���,)�����K:��̕��K�L���G?�j�v
����"�V��P�6��Nc�Q��Ӓ�)�W��vp��L���W#���#b�I����Ine"�Xx��n�?M5=��p~�����ۏf���S&l�qqz%����t�=�?��ϑ=��ӟ�U۷�E�c�� +�d�������?,'�U�I(��	w:̞����x��IUZ7�I���j�"l�|��:��7�}�����U�i���d#����
u���08����xh�$,/����(�7H�m��08���m�)��Z�2�J�Q��>�.yL��R��`�7���m�~إ�W�v���ji�I�-����ED5Mg���Z�=?���^lټ���^�n�%��$[
�����t�t>w�ܽ�92�E�П�;�'uʃ{5t5��&��h>U��6ew�go�\�]��SA\8N�=�mL��S�`up�[qO�W��R��Sd��N�h<Rd�o�w�k"�b�y�8ʫ�\�VH�C��*��Y��a����/���v��u���L�#N�W�L|  Q쀱�����g�:E�^�w�|��&/W^("�Â�|��W;��b�ѳ�A��'��<2���q���}��C�`�ۥ���SOEx��M�"ɼ��_�i�� 0sm�ă`��sx�a�I���G6�^��=�to���}��wz��GG+^�!�����J����".A�Q���R�m�n�8�-�y�.\�  ��C�U�b�k�"��]��V���m-r]�H��B��[b�̐65�ae�%���]��=|���#+���%�.��,$���3�Z?��e�i���Q��xR�ȃK#�� �GMg���f8ki}RI�ɂ�Rӎ�˸�������Gk�c�8�OH1%:���A�{�W��rt�а44,�+�2@C)^;ӓ����l>��^�j�b§�
�:�O֓=m9�5y ��U����Q��
���#�`�f�����V+f�f�r��2.X�ΪCu�<��x�7�"b��������B'C�҂弯9�?��o�Ȳ�6Pv�	�p$j��2�˓���Um[�l߼+T7.d�N�^Y��~ 2�.��Sx?��hm�7���˞�6��e���["����F@�v'LA)�Q�xp����0~�T��5�ɯ1 �m�� �V},�~�o2��1�t���E��rI*��ێ�КgY�}y���Sr �.��@w����P�� )K �,�iCj�sG�򡸭"�(؜+�.�;չf��b�S�?��I�zJ��7��3M�Eak���Y"����wϓXQo|9hRM��[��gW���d�R A�](�}z`�V�F�r����ƫ%����{4��l�Ǹ����m����b���ۤ@�;���_)*�'�N0G�m>繥���C&lώ\E~�i�6B�#fXb�g�p�w;2�5�-�.�l��T ]^��狌����O��!�M@{�[A�qw��u�{nZd5al�L{v%��Č���
_�6��D���f��K�g�uGmx��˲��CW,��R�!����:��`�p?Q�����@���B�,3��w��U��*�n�^��cM�.G � HT�Ұ�5i����3���/�gPu�3�թ�Bf{&_���r�u|AÃ���SJ&��ĵ���|Q�:��k��X�4��Z�~݌����)�h���~����gP#��@��/y������)c�"��s
���p�4=�����ƞ���~W�����T�� q�%��5�m�ϭ�,T� ��=E��g��cq�=G�
Ё��Mk-.�,�&��ѭm�Tl�Ӫ��ye�6J.�� �?Nu�WzXf�N���=��������o�_J�l�W�;Y���ii�-��]���c ��/��GmJ��j��"�!�5X����T�`bF�d��A�R �p�m�b��牋����w:D������곘�_�k�����;� �����7��.����M� RF��g����i�V=�rV
�VbY5��K�:8)B���/��Mw0��o��kiAx^��B�@{������/����T<z~���s��H/��1{'������vs_N> +�=~�v��f>m�w���>�֏���g�{����M�����Z����M!������y��gK����q�Z53��q��Ǝ�����:Ig�e^)��8ڱ����=T���f� b����;�L2�������ћ(�87�{6���&������&��<N��'< �1�����`�[[U�ɸ���YC����is�ZC+�B��~����d���x�����r��A�ϙ;��ȧ�A�me����y�oƳ��2B���RT���>%O:_l�6�;k1;M�Aڈ�t�9�赉��Y�3�VV�=u�&kT��W���5&ژ�^����M��TZ-'�Z����?k 541ԍ��U��*d)Y�)�zj�/V\c!	��s>� x�40�Va'���v+���C¯����c-&@�#Վ_<	1���&I%|����z>�z��hG-<�ѿܙ+�VD�bف/T�U�;�|E���&�xoޥ9��Zh��q�UM��Z����.qm�u8���=*����NY�L451Sc�k|�tLam��EeŢ�w(@B�S�z���ݘ���<�н�6�e���=�E��.r��)7cE�*��5��u��ށ��*+�l�{ߦ$������$Q�akE�J+կ�������+�+$O��N������˹�^
�����#pk�������?�s�;���G�I`�6� ��'2�!�׺�[n������taH>�����ه I�% ��!��5/榕��l�t0<�����Y�@�!��8�Q���Y�>l\#�2r�;#��_�\�y��F�|��?�T(�|�Jc(|"ek(�������
�&."���,dq��_�Z��������e���Σ�����d�,�&ɀ�^�F/�Aփ����j�w��$[��5���h�k�Q�5��#����>R��Y���"����D�ʼ�{�z�`��䧸��S�WB���;>3s�k����_qmT��uF��� ������4�7J�S������������{����u���W�v�q�XC0��m�1��ǵX~�3|�����폥/�ʹ���1��!CV�5�B����·UA���t���ND⃶��fR{��/�ie�/���ʰ�q"/����hKn�����v}�Ư��U|�Л3]� ط*w�5Kf{?;��@0H\Kr~�A��N��"9+�-������ߢ8������޿���O��At|pDD��f���'���.��.@r��O:��_�堳2)g�9�,�v|#�zl�2h.`�5���S����D���od�8����K~h�۟5�}j��J_ �������5�Nf��\�����_Cg��e�����N�2i?�_�_�]��Lm��Im�I0�;�f�-z����ZW[ID�(dd�'�r��� $g�߅tˇ��[���uЉB9;�^k7�
��Vi��\{�����{都�.|43~��Q��"HwA��F�*(H�ދ�( m��! -�^�ނ�@�QZ��=%����?�_w�u��Yk<9���.�~�~ߜsR0{��>]�O���*���9'W�E�U���6#�#�E �Z��y�tj��IEN�G�~�s[��?�f��Ku���{�t��o�A�"��,��D�B'y��rƉ�ݾ�ވ�j�g�U���r����#�A�����_�R�i�Fq�s����Ŭ�(�\���!r�O��ǚRW�98Lk��� ��KL�AP֔�y�}��a��\�~yQ�3t��-)�Ϟ���_42o�'��-B8u���8g�@Z��D�N~�*���qЃ�Frt�A9��R�n+�#d�����oE쓧Y8ߪ����8Fg�,��<��Skd��p�WS��r�����k�f~�	�����{+��&'�����h3��.���Hea�p_$�B!♂���rY�vS},�QD��!��i,T��:H=�nչF��U��6WG�~��H�ͱ��Vϼ"�9��YcN?���:���x �l%Dy[g��F����r�g?0#�>�ꭔ�'��1f�ӛ���j+��=̡��da˫���{�Ǉw�'!��D��5�)��Q`dY}�?��Qn���C�"���  �1��8 y��i����۸`c:�s���a���K2�:(5]����יQ�5|V�oKa|��K	u@\YZ�M���G�)�����|H�m�T_OW�mݿ�+5�Jҋ�sx�r�!�ʟ�R��u����v׼b4�5��tF��c�5F��)H�8ʪ�V�̖�U6n(���Ӹ�-ڧ~�? kU�i���b�"�2�_v��n���?��'��ʟ+���2Dq��o;�G{��)ɮ���Z���G��&Wȭ�#Pfl��*j��xO�b���G,�
Jl�)��Y6����;Q�W)�^=ao�I|i	�D���ҩX,��E!9n��g1��l�]`d�zPV��Ā��*��F���k��`A� .��%���zf>I��)V�5�ȟd7�n 
%k-��BI�#�B��fx"1Ů$J����@�c���B�mwM�	x,�qq�m��u0;��˥�N��9�2͐��YͳTV|��T��,z�\d*v y��wg�{E����׈U�D�OW����
4�/�o���@V��$�{�*FmY�r�Uv���pZJ;���#����}�jH+��U�����:.(�I�䷪o1'�3hUt$F�۷�I�3Tؖ5B�K���/b�]�g�/�B��~�|WF��)��;�`e��y�%���0iw�IĊ��� �͙���ѣ�X]�uM�IS~&�Gtw�g�N�	�Ո<vK>IL�pn��>8�z�։���"�o�UYU��S	��o��)�L�Y�W���t/}�>�=C�@`}@�� ��dv��t��s��_1+W�Re3J�>_F��8��4Q
���o	�F�O-��FFc�zF1�ԗ��x�u�݉	�SԽg��	�jE�S,�?��t	=�򕉚��fz�ߌ+7��߻ᗃ,�,hyfT��Y���,p�r*��3�]g: ���G&NIBn1�VÞp�������4��$~���rU���G-�29�{�\3�8�J5�k�a{)̊�r�^.j�.x����J���8F�tX�"���� ��$u����$�� ���I��x�+W�Ӕ���.���� z>��ܾ���<���#�
\+7'>����Ox�w�]�߼����~�B�����f����8)�S��r#3�V<{�۱R��t�KÊ�����YNn�g={��9�KUB�c���{�G�G�Y�H���ouM�� Y(�^Vڃ+�q���oZo�c��=�Q�.�jԛd)���H#$��	r�#�l�$�"{\��5*2dX�����U������|��?{�f��
`'�lN�9�r$�0�m��҅�$;�r��=��0ҺY�aeuLo��&Y1!n��)�s�W��tS��>!��	.&>~v�1��+�?P�K�Q��{�얺�u��SV3ho틍y�#-a��>��*�V���@vm��L/M+��@�Sr�Kesk307;F�W�>��������Bkc�}�����E]ԒӸ�Cg,3����v��1�q�����3+~�*�Q�{Z�]�~Yh�����w�!��&���֬�(@ղ�'VzJ�e�K@H��@_���Oֺ�Oo�e�I��avT�����(����_��WE�,�)���ԟ�v���?y]]���v�[=���7�Z����o��U�,�+Z����;~��~pk�peeWNˤ�tk�.�����8�+q�3po�����.{�J�a�v� �� �#���tWxzv�54�B98���m�"U�W\C�@��^��1/CW�i5c����S1�}����Y�	�J ���.ӿ*2��:�����s�q�х<��)�l73�,pK�p�+���c��R]�{���3���w��K[��T���k��KՊP�LMWsC=;���s}���i�tl� �&7����q�c�g����Q�l�y�g_�K�^-�������`������m��wW�k�r��e/�U7ơ|���O��S�o/w6٦���|�Q�n�飧�*��T��aq>S�,�";J�k���-�ǎp�_c ����ےd������F��"w�s��<!�!���8���W_��Ԍ�xδ6V��E��=o27s;��V��B�A����G���U��*:HSz10�H3@�nlՆa�	h]ɍ!�mک��&kooKY�|8VF`;�*��H�������%��`p�'Ǘoh��^Ff�&����`�{���[;%X�Gܒ�.:_2�^��2��u�9H`��'	�<�C]ɽw-Q��i�� �k�����+g[�B�S���Wf��	��+�8H܍I��.⣳�ՉE.6�O��;/ϕ����Z<|�{���ڢD[�/�y�>�c:ut���RǊ�����j=	g���0��X[$/�O�j ����������
�����b�$7b��4�2��ţ�X��b�v�d�z��'�j�H���T+�@�o�7��"r��H���ys��$6g���eO5S�/�a�X2ʗ�I��dU��b�,��x�b�hF�Y֞�"�K/K|	�5�K	*vb�K؈�����^����o��lx˄�_-N �}�q�	���0I3�9�S|w�n��<��뜅邻 ��e%M���jG�ṡ�[O} ��Xg������m
���(ɝ;,?`�-B򐔧�xT�� U^$oa(N@B�_���b��zCA��^%b��-������w��J��K�-� �TV
�6jƃ��)�Ȱ��fc+�Aޱ��q\��_�.�kg*$2���ܖ:q롷�(?���󀊖��E�d^��=���(��F�׺������.X���l�Z�=�t��"�5L���{�oS��+�o@��v8��X�2��DUZ��K��x����K+��j����b<)~���<-�'^f���s˝���G8H�ɟ�����֤`���`�Z���|�;�^�hF�۩k��[N�	�\Tϧ�|���yϏ��gGqdl�\���bm!�Vda� ���O�j�8@�֫����=�*�u�R̍@��y`�&�����p�*���k��`w���p�jk�>�"Sġf�@7>*[̿��a^Ü��޽Ԟ���^�o`P�t�ʊ����W�+<���1_��}�7Fy�J#� ���Ү֝�O�;�I���,�[[�؝&��ƛ���̷;�Ag��D��admQ7����&%���x�8��qL�v7Bq�n�#�H���c{�uA��0�� $"��v	�fI�[�T9�6^�:�~����~F �3��Kx�ȈDh@�)"���<���SMd}%N�kn>X����g 5}�+W����Rܜ�����v}}�����֕Sl9 	&K��O���C$�+��k�_�dv��ZP�V��}�n��Ħr���P���:�sR'�g��i= �"���J��{9�0��_�,����^qu���-��B�y��W�UX��S��� 
��6�}�~Q�TЍ�5sn0Y��07D�O�e��P��'�v�&�H��.��f���7�3x���<m�n�`�1_KE�Y@�����$�T3�mGB7����/{��u}�pMD��)����+�Z����x����!�(�:��@���Op�¿� T%ɼ��[_M��� �
LT�l]#.��6��6bv�R=�?X�|�0r��+�� b��������zS�(�k�%5H�ۡ�i�����2�C�KK�+l`�IRTT�0gt�����ػ~���ot4A���pQ��?�@h�Pcִ��[����t�b��������3cAlxF��i�l��#��B/fB��J����;H�-..FAij�ɐ�@��е�$G���-z��tj�E`n�]^x�b@�)\PPi�Ę$��x㨈z]�
!A��{�[mv|n/�3�rm&��u�����C�N䕑�g6�U��n��Cg�6ϕK���j��ޢm���o�3�-Sɡ���9Bl+�K9���2��¨�h^���*�5��V������n��0i3]
��=M'�����'!͟�)ߒ�J�j	�
o�:6���>R�� !Įnq>`{9H!Դj|o]M_�>�m-��N#YJpr~ZoD���zO1�s�g��_+=���^���qvވ�&���)�}�ͫQtp������n(V:�r#�k�_;��g�������T��S	�v�����C�4pa^/YUU����!�SnÕ���m�h��+={��+��H�C�L�3q��p7R�btX��pKt�y ��D#P�_�9��e����ˠ[��w��+�/҇5�&t��Y�농g�O�UK�Totуޘx�v�1��m��|���*{;�����RN�u5��S�LU±o���9E�Y���V��٘2,j�����1��!�1y|V!��I����z�|U[�G��7�͜;�g� Ă(���m~��t���ݾ�<ohlh4�w�ٕ	�5F�'�>�䊬�oo�3��U��ʣf��:��|"�rdׯ�	]cN�nq����3�UܲE܁q$s��׼�� �G��t���$�;�lT�1֯rZ��3�"T��S���z˙�n�7���~��)P��F*�������z!��#��C��G�z"Q�a���R]�m��:��-+#I��Kń�g�Y|9��Α>M/�\�\XR��� ��s��R�&���w􆉣��3��Q�2��@O#��-���I�-�ܫ�4�֔fsȧ�'��ax)�0`*D��x����^b��7B,�g��l��D/t��Vk~d���E�3����7X�-NUpj�o4��G�2
' OK��{��1��5�������P�}���\o�zn�z#��/JA~��a��kIto�+虚K}��Qg��݆���9��u��7�֗A��;7��7h��s�܊4azl+�Ѻ�/���f"�f�y4��hPE�@+:\Z���7k�!0X���F��$��b._U_���Y�p�JHk�����0�%ZH��Y���r1Q>�3���@�:��3Hf�.�NvHc��/O�D�8EÁv���ߗ!A�������#c����0�!�S�H�@�
�2�䢇���bE��0&s�x���_�l۽�3}���﹑7�#�c}��s������wC"�J������z��[-���A�g�`p�`��2L�>��������,�p!H�/��"�;+��-�$6`4���wD��jj��1�+�J�m]��iy^�QJ��}�c�9:�,��kjC,�2��Gn����V%���i�Í8�N�׍�;�V�B̜��T��=}:��RbފdT}������Ky2���P~� �F}b�zI⢝��b����"xiW��FmU A�����\�W�J_���-De�ˬ�+�u_���q�T8G'��M����J�։ !�K�!���FE�+���my����1�Ӆ*w!��i���,H�	�>���z���u�^�zc�Y�ż���g���n�us��ZGsWY�	m�Qm�n�hTp�a��o���wCu�Qs=y����@k!(XE9��~�ss�PHz\&/�{���m���C]T�{V	�\R-sƱ=P�'��w`5���|���y�_���B��M˛p�0��l�a��V����8�=�����M��n�De�@�Ǐ`󆧌��Oon�{�s Ȕ�r����/r��P�WCȌ����4������Ό�������QG�_��NȘ�8a�'{�v/��%P���F۞��+�0��i�}U�0��z��x�����mC�� �ăN�q8K����v����1˽���D����|��̈́K�P���w�'�% S�w��CVJݯ������7���/�+y&�����k�y�X_Uܢ?@s_� t��]�_f\u�Զ�Si��L/����q'�5>���D鍻y����@/˥1��'Ry�|9��r�α���264v�48J�ɽ�g���o�*���vns;�2�:��e���- ���x�wo�a�Ҍ�ǃ_�H��j���Xy]��o]�W�>w���z��}�07竐�6�6��]��.b8�nl��|�m�:$��6-����^�o�N��ꘌ��_!�8BL�w~��k�el���N�v����I�yE3��7��n#7�{t-�z|�ɯ��Ef����CU~�7ꣃ��� w�H��"�^l=ȇIf��Աl]#*?�t�p�5��lҘ�#�8�ߴ�9�Խ����=��� ��'�1/#�{�q=������j�K��+vt�;��À���}׼�ja�Ѐ$s؆�|��=��Ώ�_��6��sx&��Eu�ӯ�/8j^��]/�ڸUW���s�j�vz}r�6L_���q7$�-<Ȝ��s��xQ�yH3�Xܘ�ĵ*Q�y;���6����6�/�B8�1z�"Wc�YQ�k�4q����H��w@<��f������1�1�����c9�}�
��Y&�F�@�y�ck",+!G��.�&C�÷lw���K<��x�l������;�贈�V� ���-\���k�~:䎝䁈%G�P���,�N�k����ޞ�.�0���%�undf��dn]��a�Y�g`���܋���>� mb��8cl�A��~������;�o�/�&�jx�6�]�] Uj:�~�]6IL�"��9魕��M�J�Qq�.�n�*R��e�|�3u�Vi�s����K�Y!�m�D ��[u��$��7����'�.o���F��*�ް����Sޡ����	���1�����N� �W�=/8���إ$���%�
�G��4Qf�A�Q�՛B���E7�r[<���fm�.?��������{�|���IN{IgU�f��%_�d�s�jG�w�0��������S�+OA�O9q��q��G�Sϴ1�4On��7���M�j�� ��x�TJ�[���&�<G��~���
d4�3cX��� �Ȇ�z<�LUL�&b�������W�hX䖔!6��{�{T�~mÆ��>j�0����r�_�"�(���I�fO�2 �z_!@NW�}��q�_>������~��O3����y�ȷ>i���6��e�9�V��)����
n�*�h ��̍��&G��>Fa!S��/~4@��n��9G[>��/�xz���ӹa����?�1�Z�B���BzC̤,��������S@R��&ō>��]N�
��g��ٚ�j��F�tGo��*�f���j�xׄ#0+��ж�m��zȤ�V�2R��k��=X���?��X� �E�/^�{^�iqQVD�d{�?��n�����cS�U`[����RĤ�S ��TR��8�����'$(��X�"Xok���u}�D�����\�,bp��h�A����@hй�����0������]����h����Y�X�_����Ӣ@�X�rX$�x���%��c�XԓUOeL,G��-cօ��Z���(�	3Z����~�����v����V�3���@���0$(�X��_\�Z���}T��﷫��G: �a^��$���F~B�g��m`Dٌ�N[w�<?_������m"�\�q	׀>�g��z��O��3�'���
��s+�Iw����QT��P@c�� �_�}���@�h�g����|"}}|��i��0t���" ,DH�vC�ר���k���:��Æ=7ȮPle&�L�*ف
u�����RX݀��z�����β��>;�@�)�:�l��XK�������N�:gC��`1�5����
u�;c�#� �1}9�U���~h׫�6���Z��������f<����c�[g�i�0$�-,��ĵ�Ny���zR'�4�Fݎ��� Z
��\�G�$!Ɛ������-�p�� ��J1&Zz�/Vzz���ֿ�X���]T�-���/����l��sk,��D^����x�ǟ�3�K�^��N�;�x-���os�sq������g��-d���W�y�1�rY��e��	L����fW�&���!{��w7[�\QU6��]�@�^�s����ƞd#��R> 㤷Q�e�����
!�(����	�)}2g���!Q#��C�c����X\E���Q�h�������5��kR1cvc�e�� ��C͹Ț*��N�-AX�I)�cs��*�ƈ��P�Y⑪�Y�#��+��tga�j�[z�2������;oA�DM�Jc��4y���V��cJ�O�C��[ ^]���U�;���8�6GX��;�&����$�H�Ϳ�y#��b����t�e�b"�탠�P��bn�ǌ�x��X�7��yW�)��=��=�˭ixP�-�T��L�閧i�G�d���6I�67�� �o�nxb�t�����I�6FY���l,�=4';n,�`��w��_�U�+%�Bum�m�o����=�#�b��노�"j��\�)�'t����k��O�&=�f���@tq�YB_���w�K?8{�v*cF���gq�!j��eg��<���D�\�����3	|ԏ,}���r������p������k'K'Y�5�\G4�KՃFF�d�"!J�j5n_���V�]FS�����l�����>����hw�Ul����k_�Ұ!����w����)v�G�v�� ��HN����2��:�8NK\1�gU&ħ���I��L珙�#|�~`#��򄇮�θ���9$PTB���H���eU��E�jם���[ë���1W�_��^}�m�D�._H&���)�I]���݊M�`��K�J�+#d�W�^������@�ę�lժ-�u�~�iy�nk�w���W�'V�OGlW���[�5`���d牶jhO������XD�� ����;��rQÿw����MN�\����*�K�A ؽ������yF�yɮ�0�	11-��?����!�W_�����m�f�cϘ�y�r��?d��[���7O 
�C��`�_i��Ǝ:fo�*ҝմĺ^��cc�=b��J�����!��e)�t�c8w*Q��d2�HT #2i��9�zȫ̲Z�'#%C��*���ٮ��8[X�*�T�_�p!�2��^�I������ٟ���>h�����������ܵ�MJ�~���Y�㐴��Rl���H�4A*��t}a�����9�Uy��]��e��o��%�U/����vi���5����i����Y2�'��C-�S	T����\�)�A��tS}��ݱ�;�`uu���li�Ets�]��x@�j^9o�.o�D��ƪ>��,�|��,ż��'�m��&g�#g���XL���R���S��� �:��)�a���o�@�����j���6�4�R���w�;�AJ�4�@��&��6�98��E	��4��f��H�ʉ�PI��R$���W\5�ζ�	�؍U��z}D�K��ꡆX�-6s4g�b�mb���.Q�6ѷd:̵��dT��O��xɼ�,6l�-��͏�p �vM�F��a�cņ�0�����s�`�E6�ա�\�X�/�zyM��j��Ʈ�TE��ϙ��|y��+�ٮ�����1�N��F�}2�n&B�"��t��D���l1ks�Ғ�T��5
6���C$�1*0b�3���np����̋X͋{"�(��<��P�� ��e�����Uk����I�,�t35^�_��U(Y����/]ƃ�FË�y����fG�=*��8��Ƴ0���5T4�y���� l�*���X�X�]Qܽ�:,,e՟Ӓ��M7[w�	!�a(���/o����\�Y�u�x��J�i<T{aۗD`��3�DW������r�=ҕR��[\��CSyR�ƺ¬�t��+�}�Xgn��䎱�Θ����0��hv�Hh��[��ޅ�����Ǭ�;�n��Z�����R�-�М�)o{��'�)���kLJ��%]!Zx-߼�Rl�#b�#�:��}���~��Cp܆ +�д��e���fѣF�P�Pj2�^�c1a7;f�&�ی��.�F�i�yvʰS����G:s��Ꭲ�����t~���6V�M���B�Fkqp���C�����B^���E
���zwF�z�}d1�L�.�(�y��x����~�5m�?oT.95��!�D[n�"]#��.7�@"_��}�f�3n��q����X��C\�S��!�@S^G�p��@�#(��z��[�5zn�;�]ݓ��g3���Xm�9����06�~�2e�dAiX��1�w��r�Ň߳����d��<�����7ǨwW��kC�H��U�4/��ʒ^U�8�zw�:��࢛G��vI�j|߷R�x�Q��{��#̽�!.W;D��RgR*���z�e?�b8o4���5��</\�����m��k��a>9�lpw!�z�SP�Fa�n���j�a[��� 1���Qo l�˩�4V7��	P,��V�L��0Ow�f����xԏ�_��oPN��(C��bO�/�	4g6|��Qu�u�¡{l���d���CA�MFv�?�[R�<]h��H��_�\���n�8���:/%P��X[gZ�34=S�c�Q�Va�fr2w�}R�%qaOD�ce��a�n�?��`u=-˷5Rc�x�dو�L����w�	��K�����,w*=�.6��ۮ�Uo�&xb��Ʈ[QU�iO�O߬ߏ��s(f�j�mh/86(˼m9�.o����t�=��C8e��ZԱ¶�B�ٻ���eݹk�:r�wP���쀐}U]�q=��2�� �ePUB�=�,T;#���'Kץ��*ܟ����;쟕�X�>|�-���f�k�|�Y<��|*�|;�u��E�����_'��Y+g�ެ������,>�a�ݺ�{���;�y9rAw��Qd^o���n��ey>Z����h 3v���^$���{�?��W�Vǖmk�9�ʪ������L+��E��d�	�^k+��OV���d�>�~�ˣ���v���y�p(zV�6`�m������O����{�b���BZ�����T�eX�m�+9��]0��J�+�t����Pf��XY6G(u��09�+d+9Y�b�ꄍ�Yloj��a�3���:��������=��d��r�����	���%�:p#/�G��7k��U���S��ݑUO)voB���FJ��it����w�{��{�a�C���~���1����\1��p챫!��g��Q�(9��ȅ���ʬ���v��d������1k���c"�s�±���e�N���կݰq5W�-  ��QNU��jrvB��X���-���������U\�N����bY�e���}���5,��tGxu�Y��Tx�R���S� C�� -h�})����'���~��q���'��q����'ݐF޴{�?�܏�?N�8��䏓���\��B߰���ۍ�^������?�~�8�q����я�G?�~�8�q����я�G?�~����'���Kb��wuU0�����tR�׶+�O�Ҝ�t����'-/�oӇ�'䜫°Hޯ߼�uH�Th��~��%��OWj޲�_�RkP8]� t���W�YUħ+��v����z,��w����[ۨ5�_�~���߻|�����
����5��9���C�?�gK��c+���D;Hl�3����cW�;�[c�E�.<���w��+���.�#Q��P~\ $J����W�=T����D���X��Lm�����?%�1@׼`�9al��Ο[�o
.WP���i.��o�W��R�7ܟ?���25=@�q�',:}2be�V�7�}�p[�T���'Ta�B5w�C�z�tA�o��������ރ�,�'h���E�^�
�>���w����4��ݮ�A��2޷!.**J�������P�F������!�ŕ��r-�2&E�@�qG�{N�w_3�u�J� Xrξd�u3�������t?vѶ�nl�ݿY�٤ؿ����X 3���b)���1]t\��)UƓ}�
�A��p�j���OA�u��ut�����ӄE~7�2v�����oǝ��2l�j�����
�϶���X���4� i�?�]H.yc����Rkʻ���VAl2A�%f����GI'c�<�Pj��nh��G�[E4�"EUuuu��ak�������W���}?{�:;ĕW�P�<�!�"4"Gb߉��)&���s��%<�mM�87���($婉��r'$���L�Mvy�:�w����S!uMfߓ]�����*�M9��=�]
�ː���+㱌��ꎷ�^4��d��J�f�
��+L�tH-��t�20�^���8'At�hk;����q������	�a 	�<j׃���y�o_�%(~&Vk�U�kY����@@�\*	Z::�gXA�֐��z�x��S�����!�V�[O-�Pe�>�9��f�xxx�
������K	��� ���b�)F5_%�o��뉚���:}����5�wzy�i�@�;�������˷wv]W�o]�i7��W�p�:J"�o�Rr�� 3�333P�e�QLy�i�#�5&���8[���v�$t���:�P6��e�/�W��i�+VGԨ4KT�cg!��r�n�	�M�B�{�vή�����H�ґ���X@��(d�����k�uThzH2���L�����]G;nb����:�/�TT� ������\c�cs�(U3���Z5>�+PJ��W� ����a����E�n��r�Q3�e�O)D�\g~~~�<����4�ɡ+$ O��;@Ss�
\��@���~�vUA�]5���7� ��\.��B7��@��<��/{U�Q�~Z"�H3������_ ����s��tv�`��]|���!��?�/W <>svH�fr��xG���:} �j���DӜ�۾��]�j��ffJs�W�ڿ�[5~G�淀�-���PSSs}9�aߡh���ȉY ���D���PSB�\����0����g���a0�q�D��)��./(Xۄ��˚�S#@��8���Y�ͥo� ��i��%�#SG�����02�h<�0 #����q����Xg�DONø���x���%����]�=��!p �>�̖�p�c]7\*.��ߟ���9k4��9�'�XMHF��CT�@N2���@Q\���i�@��@<��~��;6P���Ls�R���%ԣ��ɭ�pӵ�W�A�6 p���B��09�M���Oi�>hb��-U%�EyI��>�f��!��ζT�3��9�c
j}�Ga�V��!�f6�x$=Х��㱫�{w��	�TKO���C&��QB�U��~Ԧ�&%-�����Cb�u۴���IN����$���É!O������V	93KK,�L���O�Q{��W4�
S�{Z�L �� x�WdA��y�WZ`oz�9���A�?x 'X[[[�|O@/<4��z�+M����g�����Th*fȲ18��P�v��A҄��my����n��z������	Oy`��e�N��in�x�wK#jiU"|ͥ����˘�L���Rz,�2�<Oʞ@r��/ W�`[�[�E~0��!/�H�F�("�9)������p�Ҡ�#�b�Ă�oY{�Z�0�}W--�����F�8|��3���c�T5A�Z�]�J،7U��}���0|���$��K�
_n��I�ﶴ�S���+�"�!11`�zW]U���_v�Z�u<�<X`.&x����cN[�s}��<
�4ʶ@�@��`N[`���չ���av���"hN䔑�@�_�ψb��`we���}�U �&|�Y�Fu�W���F�E|�=��^��ȗ�y�@8����pD>�][d�p� v��c��n�#Ǥly��`�lQ{[���
��#���7L��,-�"T�Q�g����Z� ՗�ke���&1��[@mX�<���%�6�$`8�ځ?���#�����d��@�Z��#�}_6Ix
c�%����,""��{�z����j>��- _<&:�8���Q��aa�!�@>���[QV�1�i�3m�EcژP�,3�3�x#cc��Z�u-K���$7P����'����u��m8����aB���f�2b�X���c���c��J�K��[�a#vz�0��ɖ��	���67�Z�sI X�U�A��7B+ġ0�*�2�݉�86m�Y0���Cb��|�Ɋ�.Yba��i���wIu�h#	���4ʹ�`�4�ʰ�P�/����0=�#1� @��n�E�>�e)�D8�\��)�Y�xR��Bf[FO��8S_�&����r�(EV����-�� ����#u�ڄ�S5O�f=Z׈F5�����K��7���H����ճqp�c!T�j�^N�uX)9y芐F�dM-�r.l�Na��5��iJ�4_���0&(�m:�u
5�2�����IE3��f�2�bꞽi4��zD�꾆��iH�	=��c}�
�I�^�4�ޛ.w�!�|���BzG�8���g��D�6+ ڹH��^�Jo����1�)/h�؜<q[���P4dL������n5N4�����
Cm�slQH�H {����v�kceilE/A� �������j�F0��G;��(3��j�a�8�ٙ���r�X��kC/Vk*\�AՈ�	=��G����4O"a�rv�&T?qvޚ�Sߎ�:�1,ú:����>�pqw߽� Ʈ��f]�yI�)%$FĆ���a�L533s���̯��$���@�E|c+
F0�6&�$Z]aUCID��Mڧ݇}�P�|���X��������U�Z.h���A�a���p�s)���C� ���Eh���u�$!"��QR���"
��аk�/� �!�/�v��j^"�F���JX�q��i�z]�*$_zHz&	�	��&&�H����*r#3+�R
���;>��7�c��q�C<u���˦�W�"+���t'��tͯ�3�Q+��Ht� �����+�2��,%�*�J��Vbh�:���=�bʶ����j�WZ�)f��<�e0X�v��?M�0��@�L�Л�U���(8�NT(�Z���T�e�u�����~�L��_�Q�/V~��� �gkjk��A��&��*�c8�th�J����k��<i���73$�\[N���qqo���kZ&y}�!�"��A��t�- ����/fh[o5��9��_Eb�	���X��N�!mw����E᠋x��;��Eߜ�O�iha1���W��}Ti�I�1�m���j�J���bB� �z5�huw`ѶϘ��V0��E�Uھ�W����2	�s�@l��Ʈ�v����N�=��Za���+P�a�3Qê����~&O8��S�I�Pl���4�8BǶs9�
��:�f��b�馪� ҆ݑ ��	}zBX�����~�����5�]�;؀E^V�Ÿ�,}�%�t%GC?'���BZ���n�^DD$;����H��`^�\c���ڃ��gˢ� �O}N`��.H7�Q���Pl�6@������,�F�q���dES>����⌚N��0t����oP�hL�{(g�����L�Gmg�"b�v���WWW���`%�o��q�×�GD,�!��B�<�!�k��O��}}r9yy6$h�Hj���>ͭR�_1��x�e�i�����%XM�{�5�gz�-��W�zIV�ѓߠ 	*Ӕ�VD�o�^�Q	ڏ���(��54|����Z������@�^����F�����v3�,Q���=
�.Z��={V6¶
�_�$�cF(|߷���t����t�vQ�b w\���istPp�՝��=999�n��x���
�nA�������u�H����К��O+Դ-��C���n�AY^�8�״	x����!_\_ ' C�m�}�g_ҹ}�z��d!U���Zn���^��[˕���!�Or(�
���b0b��k4d�Β�>X*"n#ו�V�7
1��YA?�ѐ�-lp<�AZek=7��ߖ,�Q��(�"1٠��Y�<v)�/5���� �͡h����{_������^�,m�9�tb����[)��[�"�R������Ό ����~��nn�@>��� �	�cCb�f���!x3=����1�����p[��:��B��>m%%o]ϊ`�� ��X�=R�h�������� �:X���$�E*J .�.��x/�Zu�t�#!&�|�Pt�aoЖ�\8�]�@�>@9�,�[��8���sh5��V��tr�JZ�I<܍t�RS�C!+%��Z�B�a����_NҺM_{�q'5�+���(	"OL�$�>M� �M� %��A��PfD��2�����(����sK
ͳ��\�QS���G۟}�S
��ǋ�􈣥G]LBB5?f�PV���p[!�U�F�֢_��q|m�!��$m�A&p��iN�m{���0СZv�}���5���2�XLF��ZB�ދ���nF��M��?$���M�Du�Š�����P~�����Id�fmT~�2F[P\��7w���@�%��E������ȉR����u)-�@�����_h�7$9+�0A������`��x�A����`�bQhW+��8<�;&TU\yuB:��b�t�f�uz��N��Ih˰$�h�f�Ä�Ā��g������L�C������;�U
�����ܭ�H���1�9��}�EX�EK�%�/ ���ښ�o�Z*��ּ �2B�g��(�� 5��hn[��)��AVD�|�Am�9`a�]�4G@�U8��cͥ���	���D����i\����W+^��*ⶀ�dorX�AK�:}��v�f�*�ס8@Y;DOu�f �2M�D$�E���R���@_���V��[( �2�1��ͩ8t2�*��3��CGN�qb�V@��K~�*qe@����HuF��XNP3Ρ����((X+�L��` <���tP�@�P �4�62��q�)'4I$R�P���}��䙲*���RrmIV�{�FB�-W�W�?�o\oV�C��
_�K��Ÿ���o���x+E��r�7�*x�'Atc��s(M�4�����n{]7���5UKg(|t�Q�_�q��t�g�+���ڈC�l�W;�e�}G^�ԼB6-������݆	\#�JcQ� ,b�A�zL2g�1ڨ5�O(���$Z�M�f�}�
�6Z+v�/I1h�\ޭ d���@?����˦�«߀6����=��/�c/ɐS��t��N/�A7�6Kbo�voĮ`���6�JKK��X�^HHIm�%"�/��@vz�{�!�xy?΢S^��Fݕ�U��pq`�@��k�ɏ�K+�qژd���8h�(?��n���R�5O�VA�_V���%M�'��u�����k���9\��r�r��c��=z�h���
 �ZPc'DW Ovz
p��'�����D ��и5��q�_�i��9�F�bP$���ï#@��o ��2e'YMO�������#�)�
�s�h���*I�|0\LMt�h_($)�����n;�.�����?V`��j(�΃�;%N� i%������� ҭ�mG�����ǽk����H���nAU՞!�2�]�-ԴDR��Faa�7<0o�þu�x��Y�R����[�c�A�ʼ��H8h��T�?����˩�0n�N�1��j�(!�ۉ���C�=E9�>��^������S�&T�A�7c���v�I��J����hh��G5
'jk���P�ǕcT2�
�#�t��Z{,��5��nՅ 9^��St�����;�ɫ�?�����jS�� lhՈH�( ˶l�XD�.(�e�n}�("�0��*�P���(2D$�a�BD���s��<���W%7��s��|�x�s�vOll�B�j�{Fz':��?��<��d�;�n���444b�+�%����S�4��I������#��K��b� 	���ÿ�1V��ד����fRՃrL�z�#͡�Z����?�o�M��!���%��q���!;���5���[+�kF���H�讋�6k�� �ʡ�Y��<����Zz�^=��	n4���2����S/�}������ݙ<�@����O��.�C��8@���'�b�) �Z�L����㣦2kz���JR�*u����c��7�V�d�d�$�*\I�P�Ɲ;���5Zx�~_���w58�¬1R5�*�Aro ���bV�*���Z�K1
p\o��U�g�����X y·zRC �Z�П;0��%onV���V������'TH'	� ܲsR'�i�8O��¾M���P����<���6~&���j���#GV����r�V�\@r670��X3��U�{{F��]'�q�npE&%W9���Em���G�n.6@2ʉ߁QTOp%��A�HQ'�3�º/b&yi��F1Z�8�c���}O��l羾��Й$����\>����B�J{�y��م�$����>m�9p�߷5Ҁ����#߷Ot�2J�J­�֨��"B��B�`���_�%|#��d��r��z�w����њ�α��X9ڴ�{`�J�vrF�w��S�]C̽�+�8���[$���߹�I�L��I����>{oi�iIf,J񕖝�m��]�ï�YkH�Y��N^ ���d� )/|�/�R�dX��St,Z�`�ĭ-i}�@���N{r��SʟlXЖn�����,� d8�/�������+���2WB�G���ca�W���U���lv��T\�� �	0U$����F��1{NG$��s���4H�3\m���XQ�v�n����$��~�2ؿ��<���`!g%�SH6DtY'�7sETɅ ?%��1ɴ	���F�1��������?|�E�䐇Ė>���b�j�m�qP�+�+	�&������qݑi��,�ͽ���
P'��Ha��w�f�;;��<<�� $�Yӵ �f�3ݳ��.{��o��E鶧�Ѝ�+�����9&�p����~�,�ـY�G֬��qf)��xtZ}>2-a���@�f+G ��͜�\b ُb��������+:F��j�p.���� 6�Nn�솵��O^��e�6�����J�
�H���w� �RsK hY�����>,e!���f��;��Vlc�:�n=�
R]�!�[H��N�Ž���J�қ�-j�$<�:����VO���S�;����E{ƒ ��Y�F�ϥY��L�z{�!�F ��S�o���=��B�!������E�����б�F�r|F�pV}�gs/d+ʊl���C��M�ʳ
	�,��@�Y�Vг-P�GCL�!�~~�c����L�)̤!�B����!� �j(d����?��-|]���1���7���+ϚnlM(��̉CmC�;:w�e/��~Mׁ0�ۮ�/unq�\����a9��6)Oh;r�H^��/��dρ�&��c��q	G�/�
-o�A��(b�'�����p�"�N1�J��nԠ]����!y��&,�z�R�Hl�&���V�<1Lx%y����Pk��ZrL��wb�oz��c8�ϊ	�>ޗ�!mF���Ml��`7���'B8����lvf݈�{��Iq/`l[k�cNH{f��u��_�'�8 �;�Ly��D{�\���9Ґ�e塭5ڞF�<2A.����7�Ԡ��3-i$��[¿�	��YV�/���@������A������ui��ّ;��g��D�Mƍ����\�����c�Ϲ��߶�P�?y��˴�.�1S��<��F���5���W�^mV̚Odw����2-Q��p�Ih^Bd^�$���$�~�"�Y)5ѓ:t�h1�*��H�p�mQ�n�}@�v&�Չ�jtd>&�,!3�z�apH@P�F$i'6�e�@�GogH����I�;�`qz��y=]2b��fa݁��~�$����n��P`V����J:j��Ǵ�nbP��|�����L�@C}�e�DV��קf�k�!"�y2�՛K�u��0^/a0T%y�7��:@fu^w�
�.�Y�������Nu)�>B�;l�V��t<�B�K�3!��/II� �].�8�.�FA���N+��&�#�\I�~�"���H9G��h���#�/�qu�fu�ܨ�#/�kz8:U���)�L"��"�-��=M14G��e�p���CU���Uu~�H�-�Ԭ���r�	GEM#���#8G}� �k�����'/�|1s���h��r��*�$��	��(���%|q3�9V�{�x��{"��ɔ6�}����<4��T�F��B�hK�������ȏ�Ν���Auܷ����j��ޓm!�$=���^�'{�3�-��;q���G�p��W������npϢ���Vn�m+�B���hiS$ϛT�v(���R��!M}iT��*�8�-��IC���X�[��W��J�f`�9����ʊ�BҍfQ#�0�K��2[KK�4�)m�੯'�s��3�ι�����1n���ҩ�sK�,��X�}n�؍|��x�<�.�g�"ZD�p��А�Վ�ېJȧ������h���c��e� ��{ ��*A�9��/?�����`-.W�
#�}
s\�m������1�36�(��	��=����w�3�L��)����<?��d�bʙtY
��!�UC:����f�L�̙��0J�U<��V$㝈Ŭ�;���%H��@�;#B=+����+U�&��%�{Z��n`d,�R/��g��	b�=hҽ��ݰ��тS�������(�I�R=�6_�MJ61����Ȱvp�z�l@l;~ �WX�Y�'����`���տ}�puu��a��<���ei)�G��P��,������!��G�PDd)��[�r\b�>j�)�H(]9���.��֚�_J>og���]�*=����s�vl�+t�[E����ܛT���K��4@���I�PJ��|�g��#��Bm�����b����+��zޭ%k�WY{@4���1t�Ԡ����Xxh��|CC騄���!��<A6/u�ȑVAѳ]���b��sRj!�C��Y��nɀ�`�hY�Li����Y�$p�<��5B�_HO� Z���?����u����ai���Ą��� �EzRgv	�5k����|0�E��������t�8�0v�!6T{�uv�x���~T_(��v����`�VB�|�3��j�aO���� �]0 %_!*0-��D��c7$���
�B��, <߂ceRb�3Tv,�J�����.ZE0-����"��1����#��W!��]���~���<�R��*�LA�i�_��-=.Eۂ:��R����h}�}td;����d�I��>��	������[��Y�g�b��k1)m*���i�<ǭ�'*0��b���Tz��&��Y"m�k�d��uMl?N�J?�b�����{�r��Ԯ�\��������Vm+S��[V:h/���Hl�C�Dt�
+��K��Il����N �6��$��h
x��=1�*d��/鲣�P=#�%���4ߴ'��%2����V�Ỏ�ДY"���>�����"��v���LJ�\;	2�!_�j���+��s���9�Im�L?l�Z��I7o��?~�U4z�.SCz�r�\<kzd���#�A�,�F��9���JMM�����t����o3w��X#i���Ga[�?zZ�V̾�n{��s��DD1��K��@ ��<q~�������V_�v��^㤰���fy��k����u�������'֕$���c�ͷ���g�
\��ܟ����^BL�$�.ax2{)^��#7'��-hr�ߵk�J��|�z�!b=�ʊ������D�A�`�z -��Y��\$k�ų�~��Lw�$�"f:�4�U/ͿO��JDW�e���'L{��$$�,==i��jǩ~� �a�2F�m�_����=-�y��|��Ӌ��o�G
U����P�C@จ��o<����U��[y�U|,N`D&k�Q�е�̢�&��̓ˡ�����{ɭkZ� ��w��%���P�S�l��h�����\|�����1J`��C�o���޽��^]�����LAC�&$�+�7�����;��԰�As"���=3�"��U�"�/"�"3E�"S���B�A���Z4��KT"cPź�_#�Z�Y���C�p�L�wӽ#S@K�Τ��N��� W�P[7���!�������Z��C_텍�g�J �*�Ny"wЊ~��>&p�b��M��[y��Y���S�Y=o�zk?�3��������j)��ﳤ{�T�v<|��Hs#�A��#=��cd�Kn{���wĢ����aYkc����*)3;az��3��N�&��V���3�g�(���R�DY�<�j�J��ˤ���̍�F�ƭ0,S���X���A[����Y�m�v����ۧꨓbm2mW^s~��0�ۄ���`C��|���9�}��'�})�|`�P�!)��v��,8[�s�W���\�QF9�P��Bx
�!�^�.�XI�K�����q���I`�����_@5�L/R�ۭP�4���--���CJyE��>Q����#G']�:ZEc}���8���1�;�p�6�'r�JP ��$��:4�y�r�1���fLS}}`/E1�A���AA^?:: �y���^��a`����ɞ2�w����h�؀78յs�����팘^��2n�^��$i{��^A�������A�qY�]���6L"|��K���G�OS���lے��#5XNl5��޽{�b�x��&�Ǝ���w���]�X�_��R�D��$=��g���"��$r�[Q���z�K�jMK��	e��q�Y2�9o�<{O<��"�=K1�H�����E�e"?���[����٤�S%
�d:�S1�Od^�x�a(��U�ۖNOYEf��!jc����Rm�"d�1�o*�@^�uH�~��i�<�j���7�m������39f��Q7B���9�<F�5ՙ?S��2N�O�b�5onwf�C�,QoݫH�!�0�l��i�ɣ�}ן�z����lTd� �?ծ��D�������υҷ|S���}Ə !}�p��D���vi@oS�~��)� (c�~T"b�?�	�7mڴb���bF��e=P�bW~�e�zm�����Bz��(l�@��l,���H��l608S`�V�����4�D�7�0����C�d����K�����C;)��%;�����ߥ����\.���*��u&�J$�԰��'����_0��sK�~;Cq��f�?Կ�������23Ť�ِ���]�ic����󕞹@d�%�RO$���3������=-��'�b����j˨�(������"|^����|���-���y�砯<+�:&�j�*��������������3^M�'�If!ũ�~�!=��KC�$��xUm�VL���!A������b0i´؃���[B(%� ~�Xob#�Q�u��̩���,"fB�se��4������&�
c�^���=딏����W'�_�d�P�7�evD��N��<����EGH��Ԏ�~O��i�rAt��'�&��x`~c�{t7~��z�3��~�|T�.k?D��7��n�r����g�crp�!H����-�I-�[ๆ_����7��z? �\t��xlHu�h65!K��<E�_yz�#�^�ٴ����"�P'�h��,-U�>��a�~A`βr�txl�	�~�4@����F/���$��]�Ł�ԡqb�������({"� ?<g4�S|���¼A偅�����qu7�N���S�:�Ȝ���)�х�~�X巷���sfe�^�c���?���l�����˭D7l/�쎚�d�_.��ߩ�s}sV0���tj�P�)jz-��������~ ��.��A�]�R]z�\g��+] ���p�<��|
B��]��.��s����SdG���'U��r~���"ks�%����A/Ÿ����<H��]��4}��:������
��5��8CZ���3p�r�?���tK~f���EO�o���Ȫ��-��}�%���ƻ��ԺsC<����Θ��'����I+o��1�qo�2��"�.�ųH�[<��	,�8N��K����!ĉ�֏����v�8��(�����#Ky`d�����u�*ю�������s�q�� XI����p=�&f1�cG�(��*�5�e�����r�ܒy@oUѦ�#�Q�>����BQM�����FԶ,˺3��N_�O/ ֔���ݑY,-)\�hJ��rj��=,�'�ߎ�$`Y���o�_�>߬D�:��*$a+�?�E����$_.�1�v-`0�V�����Tk���xv|H�`N�n�\�^̑�s����%��w!tB]5�������f��l@�b~'����ru��ˆ�v���2���C����3Z���ѥ�u��>��է�r '����-�b�)]&��`��:�xS�.l8�y�T��w#��1����g����ͅ)gMA3Q�a�fQ�{�P����zg��6���� ��l� ����h1�N8pqp�����a�杻v=�c�.���a#��w˻�SR���ּNM� 6�d��"�}ҟ[;�-�V%<�<?HsL�5�0�?tǺӝw \(������G�r	#���ϟFcŨZ���e�-U=C�H��Nk��.�e�7u�̳C+�����u��������5�=���L�Ѻ�X���#G��	A�۠�xBU]����1�>M��<�Q(z��$"ڱ1|X8Zo���]��ps�MT����9z\�v-d9�А�N1h�R�	�P����<J���q�=�
�N����b{�%��!ێHKg��+��͛���f%������i|
R7{�����aZ���Di>W]�9�:��M��P�����Ԅ�ށ杮KF�]f�7�B��5�,��'ϋ��ģ\Jއt�L:��y�f�\�nQnn��2b�|����B��J4�c��p??�V��o/���hJ<�ߨ��wl d�nD3zb��x�֭[Co,�4���K44?Ɂ��0�D�{������S�\�ʯ��QA\�YHrU�[OX����~"�p��f���3��v_UoMT���� ��l���f55�Z��(��l�cJ��g�）�H����Kb ��*�}�������-|]�KI�&k�^�P(��*�������mC�SW(U���k� ���7�0���/@�KDv?u_ ��@�PtM��f��a�Y.Z�(��k/P�����Ϡ��p�9��I�9bJ��|�Z���l��	��4���scM�RH%��$�)0X�0�㲗=�gG�BG顤U�ӝ��h��N�%F�B�)��j�n���;f������`�ɬ�j:�;ml�w��򩻵��
󚆫+**4�lb�����T c�a#�A}7�r�0�͖�C.�Yw�ޭI,N�w����o���^|���?�V��HuA�iUY�'�6iū$���(��Y��Ь[]�:�ԋ�0�5�k�P����C�	�_��T	ވ��S��o�����Ϗ��8���2����tde���@WU��1-�cs�D��}��z�Λߡ�)9�%�71Z����"!�Y"��d/�V��]Ҕs��!w�<��_�1n�����e �\!m��QȨ��[!��	�	�Ro�>|�1�V�r|���ǌ�5����Ϛ�dee�!nQ8�Qq��0&S�-��e��D��n�52����l)��/��b��2V�l��P�M�C�����9[?/��X,^�Ou�c�{ޔވm<�޶��C�p%v��Jݞ�E�n����xb�VH���'o��tp��@���ng�|���.���n�أ�7��x ��x�-�����k���UN:Q����� ��7���R[I�1@Ԗ=��e�!�Re\�]
|s�ʃz��j��ё��ųS��4�R3�:�[-�(t�Z$v �����k�.Z�J���%��.��j���W�L2��Ԥ97n�:@�$�����Z�f��`qQ>����
�a<�iI��.�����~T�(y��� ��*��߹<����㍘��/�Txм掠�� "�)ڤ�x8���1B5�Zw���ˠ��Q���r����h�S�'v�$Y��W��\PP0��;x����2��E5����A}|����@�� ������u�qn��\<�)�a?Gy��c �t]��Q�D�l�e�-�~��rW�NޡE+�Ju���`�;����!�Y5��t;ā)XUB��Gr���%pÉ�#� �X�YoHߡ��S<��')�e4Y諌�������CS��duc,mx�;j�9r�#)�%���B��eD~u6]<�ooB[yV?A[�(s����� ��o�!�;v@8����`yRrl�;e�E�Z�8�f���P�C"}h�#;D��s?Fk,Y����w+66v�*��a��@CC�	�Ԡ/1-���UU�%�F\8�*�hS+��i�K�����������69ʫ�
<��A ߉2���6m�8��=���9�bJ3��&��xъ��@���Esk^"��Q9g3X�{rݖ0�ȘU�u�I�V̘6�(W�6�S��?-�٤ &����e�#2�#;��u��.ʮ U끠�)7c��/����}����������4����Ё�b���a�a'�vݘ��g���aa�(���tv�8�(�BT����0��D�w&������mp�����}ׄ�����P狁n��6V�ǜ�#�m�h��1���C���:㍑����x"����H�5�ږTP�9�ʸiݙ����#h <R)cz5a�����{b��.Yz�oò����z:F�LJ��7�Y�q'1�5h/�)rI�%����ץE�B��hMݩ��i<��6w��Yu$?m�����T���ߤF�3]d�D'��{���>��EM�P>Z��q!T�_�ñ�̊�<QT�*S�1�@���F��w� �o��2e�y���:
f6��ai5C���՞)X����H%H��|��3�mb|,ެ$	�\��4�A<���2�ʠ��Ϟ=���VhİO�=��w@L��?�+�m��D��,������H"��ug�I�5�J�v����CG�U�P���V��u��(k㯮!�Ɖ~�r�?!�Ӥ�m�b�����]�?ae��2�)��C��|��`b��xOHּp��N]�z�Çjݒ��3�@+�n�p���;;ZP�Wz��z�ׂ�O�d��\��(u?�˛)u�����첔�
X�������}f�
��v�.D�2B�_8CE"Qfy�'�Њ�ֶ�=򠪫�j!k�ۍ=�q{�(�*]%�(6ԡ=���{�c}���L�$�����&��ai��Ό���(�e}��zȝ��A��D}la
B�A��[A�%]FK��aЛ�i|�?�U�W�u�þc����A��:uDx'�cj�+�A�tY$�V��CFffx0XjՖr\�7�"䷌��%S��3#�#P�#�m����mN2�Tϸ�f(����g�m���L�1/SU+z{)*�7;]q]]�6hmI%���vG*T/���ˡ�K���H�+)#mV�5=m��Ѩ�H��nUi�l��ٌ���P�:֚y���IrCÄ�v�Z�SMAC2��Ua'�K2LJ, �ǉ�_CI�ɯ�z��:��:TmQ���J��BE�ж���iGQs��mݛ�Q��դm���(k�#��{��ŭ������j-�c�T뷸�U�_dRRK�{3�u�/�鮯)���6��ߒ�sH�[�x�ྜྷ��맮Xg�@����o��g+!�y���uG-
�>�!�1�K�%j��e�"�k o�'Q3��{��y��G�?"�����oZ�v�
��Ɛ�� ��JMK��^�7o^�9PzV�[���?\9,�����*����L?���פa��gcT(��g�V�׼�C�����.Doo��u��ug,]G�z�0��Z#��Ep��'��3aX���`���i�P!:�BF���:��(��jpʺs���̀��F1UH,�ynn�~֕	ԁ��Pw��*h�Y��16�H$�2z��R��c��S]N>���CI���^�q�����^�nC4G�lw-���1}���t�=���s�"�,9C���� ��5��<]6�UFk��,=iz�3�.���5ϵ+��
�U�6H)B���,�0�� ��EwI�Y�toB�9!}P�D�Q���U�އ�q܁)}E���RKgM���v`�؁s(B�}��W�E��*x����*�V�� ��1c��D��Cew^�;v��c$+ӓp]��E�x�4$��H���t+E���UZ�����"��ٿ%�w��N>Za��5 �H!����tz�II)pQ��΂�������U�?|-��Vs�0�Г�k_�X׆ҥ��:P��eR�y�h��Ћ�\�������Oz�|���?O��YJO�*�e����C+��r���<y�{EdO��a߲]�w����9)ݪ�� Wa�� ڒ�����3h��(���w��{�m���E۷2�ēP�v|�%�9����#Z}p�B(������7��f6m�QәF��R���N��N]�쨾lV�	~�r�r���T�0�������@t>��hŇ)7fݾ=<b
B��;i/݋��6�1�ڕ���߇Xw�-@c0���aF�x�V�����NO.굄RJͼf������Jn�����q����W�?^���jn}�GfHp�������@��wіn̬`�}���C������s��U��S�;�l��JW�j�i;�m�w/��55�Ӳ�2OpF�kb+g���4�6�-�V[�G��3�q���ÉG�Y��Y7��8�[�cI�>��H�v5��ܜ��
�<n��fp�ԝ�98�8ȝ݀O���d�O<>}�I�~�]���|�II(�k��6/7�?9�����MvM���@��}~���p�O���q�Ol7�%� �^;��S@CT^�:Q�
��7�\O�޷a4	�]GP~σ�ל.kP��W�~������Kb�"���6::ڳ<�=i��P���[D��j̄@��L��i�$7�Κx����V�,J;U�Z�(��!PVD	�w7M܂��xt
�ߘ�4X�6"�S_�})�b��5��J��J �*���b�R����)����T��ž�|�W�u��R��Z8k��H��WU���&MT���C+,����n��j�G/l4_�5��J�����2�	Ɣ�ָ��t�7��G �����ne려Zĸ~���!�L�F����������e&%��Etls5-(蕁��L�mڦM�R��',E��5�0Z��ɩ�?�=�u��2n �j���A]��E!��G�]~Yv~�������~wwwC�Gmj�T(�`���dH�b-
��ֈ��)�EB��}n�y�[��Z�h/�;��͘Z�6�;��:�+z
��RfۮP�P�_�^,c�A�
x��*�����xA�k,) ��E���>�m��e��S�Om�82V�����������F���0��{�w� -'l��ԉŅ��?�.%-�T�{�{S���GވBԍ��Z<��LJ�*�>vuJr)�x�/���ݻ`V���(I������|
��6wdk$I�zVƛ㬯"'gPvo	�N>��:�xiii�A�>A��:QX��X�h���d�4`Q���EY<&ވ#�})��0�L��؉�_�Q5�o3�IwI�h��͘�(à{P�z�uT2�Y/^С�I/�c�;�w�^��G��T_(K�%��{c��?�0��_W�^(~��A�����%�q*G��E�ˁ/���52af�C��9�����e؟"|�Ỿ�YؑJ#|,8W������'��ms-x�8$��r귁h�/Y����P����S��F �y$��OEn/�VV[����#��IC`����d&ɇf@9��H�~��h�öQۮ���΁R5�]b�3%��ۦ�c�ju^��Tߣ����]s}r��V|�䖋�:R��1�ut�9Ʀ���(uG<܋�m��th��:^@�:��b����~S���U>�܂c�s��Ռ0&n#��*�-�15(q������� Ӓ^<��U�I�)z�/�9�x�}rCSS�zEg�+CBD�ƩM�]�z5�ڵ`���u�
�o��Yˀ�j'�"�=ɳh�_{Y�G&�Ώg�v�♧]5v?i����q����[�Qs�{��ʶ��E������;ߧr����"�Î{�ά������_fݢ3���_�j�����]�q`��}Ng��+�/�R��<���ƒ{_��h5��j���8}.d5�(P�u����r��8冎k��na�0���s@��`;F%�ŅI[�4�eH/�����s�D�75@C�\$�3Z��T�<r��0,��Ra�fq�}�X,�d�:��6�U��|Ap�1� ڠi���!M�x�0�o��#�¨�.��}����5h��:F�-�{13��d�/$��By%�/�P�rL���E��;�,; ,B_��s��2�.0�	��a�	M�q��Dq�z(D�=a�Q�60)���&��]�Z����=���]��Dw���}\#��������+�j}C�?ѳX����C����������u/�{��:t@hܜ��;0��Q�^���*��W=��贺1>J�9�Ժ��0�Q<Hd���3�OŻ}�U!99�<����('JU���{|||���e!���a����J�)/x:mI��I�z\���9ja�� O�P����gόc-��2�QV���o�)�]?�݉�V=���M�5 1u���L	#�Ip�$�� �8� k��O7����ar���@��OBnS�#��8W5-�ka���a��X��T\�,���l�blw3�0���)��:|��,����]�z}S(��ߢ�5Ƽq�[�9������(�e}����)�g������}QSq���{n9��ȸ��(�@ʯ���"��|�C�71�V	�`���7�?�m�\^��S$��5|b-�Fޜ�z��3�������| ����WGa��d�7v��"�,ժ����Ng�fv@�x��%�6݌����
v��e�C!~Ѡ�	e�# �Bk�9'��D��vI�����
*rp����`d��7Gu�P�d���=euHS\���N:�b��g�61�LJ��X�"�"d�)!YK�>.���Q8۬]̶Ԯ�T7����K�+��)��0�C(��r����EЧ���6S+0B�N�Ѧ��K� k2dl���������*���'��a�Wa�/W�}���R]���u`�/F� )��O�r^8����gڢ����f5��e(@B'�x	v(�Λڟ����ݵ6�*V_�?8x���T0���yi�����o��
��y���y��+;��G/�v�:�L��k�Ǣ��������{ø�8��\�����@�����k`������'������*�Er�w���՗K	 S����sZ��E�rsv�6B��!�"��C+55�(�|�L�(���o���-��w��r%^��2�F��_��4�K��@+�c8r���|z�]_-ڴH����Xͳ8�_�o"�����Q��20�7��g��w��2�F�SN��0������nb�T��'Х����a�y�j��V�u['�r%�\n��P>��d�� '����#L��Cv��4ۣP��Po퀝�����u8��-���Ŀ0'��47��y�r(��6�z׮�-�R��j�dqMP�L��t���*�=˞�(��t����1f%���샵�Vk �S�h��eee/C�����VP�Xa
0D��8����vΐ��c�o��S��u�j��r�@�?>�T��O����#����7X���ao9螺?�V�J�DO�c(�7��W�S�̀�ĉ٦N�F��ns]����6��d�Yǂa��������%��'����+���R�D����$G$�WX=��wW���)P'!��N�/�}؀J�����E ƒ).�ʆLo�&�.�
���}�ԗŹ�/�7�=�OL/W���R�5'�������.�u)U�� �zv��17�/���ۦSǓh�?Kr3!�籟��~���wa��"�d�Z��6�7��}�;�1*������|3[���ޖ��S�'�LA�����9Cl������T���v�L�)n���#��v��O�:]f
���6�E�}�>lt�b���y^%B̒����\�e#��c�Ae��������\]T�H�_�����[��ݻs֮I��ܦQyMŻѯ�p�r��}�	GJO�1j�窤��
��"�����������+���̢��6aڌ�+�J��>�h�H��ԗWoڴis��3��~>P��0C(.�O��F܍Rbr����%ɚ>��غ��!�[kS�8��%-��u,V����X�.����8�)8�ywC�e�e�� �GP.��;T_ҵ��-�K���6�O�M��S��c�p ��|��q]��� D���}��9�]R~!�e]�͚������m�q��&[�?:��� PK   .{�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   .{�X�r�44  /4  /   images/863c2d63-52da-45ba-83bb-7a6a6689309e.png/4�ˉPNG

   IHDR   d   9   ��}   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  3�IDATx��|x�Օ�;3��h�43Ҍz��fY���c�M36���ؔl��4H�f7�P�d��n
� I���t�1w�d˶���h�M��s�X6��g�?��Y3_��=�=��I�w�)��p&�:��ˏ`(
�$��z�e���}��Qz`�NP��G��ѵ
�A�>�r�J�]�g�w�8P�c����1dG�R��\x��w�%u���F'��
Y��"�g|�F%��]wB��DE�n_}cN1�O;���_�|/<B�(TJ9��i�°�PI
qO����nY^�k�t�5��~�g�svf4�L^\(�s����?�*E}�Q�@������@TäS�D���Q]h��5>�9�?�!4���ͫ�i�<��_^ZJP���:Ep�5ӽ~��d��	�`�l+�1~7~:��P ��.��S�s��9lǕs�q�e%s���W��p�!gM��?� ]�ii!V�Y�P[�����nTv�
�|/&��e��}e��جor�C�;�*��e`!ir7/)ſ�8��&�}O�| p�T�Z���OGj �t���*|���P�T[I�!mΙ������	�� qӹ�d��G�Ɠ%֗f�+j��{����Y���ǭc�[a��^>&T����=E��yXO!jw�@�$��x�eȕj��t� jܯ���JFU؂������5���(��A�'DcC�N�y�)�s��!��	�|�4FEY�EJ�
b+�;��+�R�}њ�f�8��d����̪ʻ�-�����RuCI����|�`/$=������$�������/���d۬�#+�s����b�@䐻F���eѿ�A�H(����-L�gD��n��B��$�2�
5"����h��`k��������y�2�����9OX�Iw\S�T�cʛC
t��ARi�7��J��j1�<��L��d5d��g��8ֲ�9r�[D�5�)�����I<_�рeF�u%\.7�V��"b��#V4h�Ȳe�
�U+I�!Dt���9�`�'L1���c|݂"

��'�H��/�/#�<E�7�?G��$�(���N$B�TF�v�� b'/^�X8 ��HR4�<m��'�ͦqER ��a|�6�t���+�V��'�|f�p@�A�����FQ`FA�
u
���E>��߻�o��I������'�3����y~&Ǣ�����������wl9%Y:8GZ0�҇y�@-
��)F�>�B���Bԯ��XF���</-<gƖ1N#�a��\,�E�4�	�}h�zI�{�Z)�5�k�E�N��t�] 8�`xŲ%�<�E�F�s�è���B����rݺu8�x/������3�(	��ʙ�	������H�y�#�����	�pP-���r�Q���N�ؠ���z㸰&��S���8��C�D��+�?���d�x���� kw���f��x�|H��a��p�c�c�ܹP*���Q�Ø]w�uhok���?MI�����|�y{N�v�oc��koEn�py��W�X�,py�E�yQ��	�Rꠁ���M�[�����uf�On��bƏ|j�����
��Dq",ΚTUU��/���3����,(��*d"��(�'5Q���o�j_����VA�i� ^;ЙB��oFTE�J-�;��N;�dR +_"��oqd������<o���TZ��M�ҍ_��70��;|^/)�F�[̄�hƌx�c����� �zb��Ā��������tĲ����3v��e���$:yhҋy�X֒���3�*�;q�kB,)`#�l�zh?�C��S���v�ۅ�'Q3�6��$��`�*�/]������V�P�)�!�I������7�
"ߨ��%s֩��Q`R����1dg(��Ŋ�w���c�2g�qiES�	\��2�U�f��#�i\r�#N%�AW+'A���N�kQj��c������R� ~?N;���
�]N�ƭ���>�˖.�/<�+K�bW��`8E��'�;Z�q��ƪ����� �Z)f��J<P��)����b2,��.�ß;�����Bzz:�~�pOl���P0�)��JE�M!�lAwg;*�J�Ν��m�aL���)��ͺ|�`_F��L��}>dR�(2)1�bA�ݶ ܁(����=�"/����IԖv�l�$��F�}^�fc�W��k�4p�4�����j�~����7��C����e�F������7�)�����E��+(��� T*5V^�
o��9�W�o�N�+�g%s�}��ВW�)��Z��#�t�)�����ra�`���l޼�BS�ш8��`���Ğ���}>/LYYE^~��RҚ>����.��t�p�4L�O�w,��gqe�\$�bW�OI]Ϙ��,Zz�"���ꊳ�td���:��o����q�P\��$�Ŭ*
Kv6�/[NZ�౱�ͻd�pYa�S��%e�O4��Ks.*)E���8É{�P����6~�"�^$�G;�Dn�J!�}I CȜ�8B�$;{���&�&�_Y9C���3g09a`�@l���*��Ҡ�����I�� �`�sOa.œ���c|��W��'O`�(���B@"?�K��bl2_Y}=.��F�Vzm� �O֓I��K�_7] 4���b!�����t�l�.�I����F#N="<+���MX�d)��3�>��f�8��2��G�h|@�N WGrM:�`3v�'B}1j�
	2��$Ԓ��L'3!��� |)�ϲ�J������s
Z�����r�r{J�����Ja�,�X�z�DB&C\�9ز�)A�c�)�� ]&�R!�t�1�2����%�����1��\���n,�d�V`��BPȂz�X����[��;7�2�3�s�򑝓Y�D"fx<n"5iB錦L��*���"�"���cG�,�b���فI
i�S��,�H,�1��ntQ�����3�U4h�V)ā�cx
^�.��#��jo���G㑏�P��j�zb>��#3�(|p��������=����:a���hAqf�e��y|��b�윂�,7���r�%M+�DNmԋ����Zw'�&3���0����
�0�#j|iy�Р{Њ̾w�Xq-�am��1-N�*�I�0�b��o+)V�&1�y���dJ��=���3���B(�yy+���̹��IW ��Z��cd� 	%��1I!��:`���WT��wv����^�.h��f��i����Oz{z��W�rr]�6�$��W��KN�'	I��V��].�8�9�.��d	m`S�)�$�AZO4�qU����/���d
1I�͚�P�D	&۔��tp���Cم[e��D}��<�^?,ᣨ^����{��9�I��)���i1k�uDj硁�x+��@�l�#9B #�ᘪDAQ� �c{�V3�2�bLF�R")<��]�^`���M��I�՞1��c ��K�2ݗ��i}�P���Qld �;z���Ѩ_8�i�j՜"QYe�ӓy1K8���щ��V̞33f?��q �H��&?��^�T��w�!��B�ϊ��P���gѮ9���	���n"z%T� �nC��N_'�F���ï4���B��@L�?f4�6�|%��~�������K�!Դ��U��O�j݃�0i��/��ȋ��~,߳�-6���XT8>�������X��*���`o��hr��͗����F���Yp^����W��?��y�l���C��2r�Z��N����L�%�����8�2��3M���`�P��?��$���l61褿���s.q��QR;?^b�3���pS���{�bG�����m;�}��~��<`PZC�Ϙ��4���Q�{�cO"2�K�6mCh�����|ț�Z�gя_���:���i�-0�y	ƌ��\�C��_�dMza��=�v��Di�,����
��I�OL3-#K0���r��j�gj�0�,���e��qqɣ�V��V��^w窪����2
�,!QzP���N��+$�>}u���L�b�\H�y�<�,b²��Q1kQb��Ufx�J�p��*����B}!�w8Ѝ�7P����B�� ���<�
1��}�a���Ԏ7���	dK`n�QSoB^4�!ˏ����z�gI�ggg'$r����'6�Y����]�Y��%���'�Y�����5�a�������I?��>Dy1���W���_�1�Y����0�)4�K�@m�	wL �(c�XRYY)266&2��µ�<
l�FL��	-�ɐH=>�����,�b���z�������潐gW@Qs9����- ���F��z��߃�������S�*�AQ�Q� "�g�Vy	
[O�zC.~�-J|e����"r^2�JX�S����.�e�21����5cnN��Y$��$
�X^��P~��рk��#��./�9�cH�L4.�&�_�4���Ξm�L4�eegB�����tZaI������
��k��F���<�e��&�͛�3T�.�J�Qkb#-����d*�]yV=|������~�4k6���5��5��h:�	J�(��� �7���0��� -�5�DT�Yfʧ�����t
ϗ)���D�ٳ¥�C�[[�-@a�c�`q��������,��cL�6,�2o�(�m�w\5�^����V��nBiuV�rQR�AA��l���(۲e��G�5�&w"�I��~vi����j���E��'~��X�<(c}�~��,*J����ɼ
O6�qut��3Q��Z����.-��W�&��@oKZ�!BVu@��wV]w#��0�4�BL�%\�P��]�h��G����0���d�1���z
˫�;�����3�:0��=P�����v>j�t�Uu�#��ijlZY#�b�2Aң䛴�������d���@�� (S�:G�o�+d�!t=��S�#(��:0d�O4V����dYs_���.,�n���߁i�0�>��4z���4HcMV�.@��
�nW��u��,��=���)�j���,�p�}��}x��ڬU���++xm�(�Τ���_�(0{��[pb(@�	A
Pޕ]�1��9�XW� |�p�_�\��()d싲��0Ҫ9%x�O �$-v��i2S0�+Ri҄���Bi���'1d����Px�W��H ���r9K�^wH������h�L)�$����+1m�vm	s�A
�u�S#��;���`��	��7���k\)����BSh��'O@`3%V�8m$�J&X�ܢΥ����Ʌ@�\M�EE	$���GCI�y��� <h�$�E�E����\� �(S�N54v�)��y�9����d�=����]��u�������²|,ep��Q.� �4J11����H�"�q���^�7�	��l��0$�-��#&���$ֺ��y�;:�0Y!$u�"ˁSD��[8JYLd���I)"���9;�M���b)�?&���a�U���L@(&�i.r����{OS.%�:适\$1 ��sd��')�GMTB#geTa�����_\��>ڇvM9ʗ�"��s��	غې9zO=}
�s0�܂o�d+���l!�L3���1؍QF!�_9f�z�|A����K�|k&�Q��+*��k���d���v�-�>�F��- ���9��47����w9+Qu��x?u��Z��2(���OI������L� K,|E�1r�
��T0�߼�(ܦ�ۗ(�%��"�|��J��q�z%�~�?؊�<tV]��.�mw=A�Cn���"^��|��GnENa6��V�^�o���6���h�Љ#��pO��v�S�_T�4E<��!�M�Hq�D�~�ɂ��jQ	�(��<��=6���K�%4\�W�_�o~�q	e�s��"�փvm)�0�S�<D$ȉus�닽���C�m9K���o��7���^)V8�HnJ�G㫎ܻ �������Rt�$#.C�$���P0w!����	lcƚ1����T�YJ(�Hó~s�)V���=�W�:��5uH/�F^Zv�I	��QS���	'�X�#|���2�������47�c'�(��/QX������J�t\������i�$|5���t((�����;�S�J�K7��軐�~�r�	[�nA��p"m��c~���m���2D�>��;�Цù�E4X�bK�
G�LB4A�D=m���Q\.����Cޥk��m�J��^�j���~UC�Ҹ���˩�����?z7߸>��y�k0��	B�c�h�)ܩ��R,��e����m)�Y8Ϲ̅�+I�\�R|�`/�񲼌�����C�/�݆��mDp߳Ȣd1�e�1�B��|ь,�y$�;ȳA=�XZ�ZD��4��?����bW��8>�	Od��I�.��D�'5	.�F�U��W}N*�.�JMZ�
�ysp�=O�'�[_ߏ�;B��P/d Vk��ɿ�^�;Z����H��EE�y���2^4���$A�S�YX��.�p�,"ީ��
������U��>WP��n�
'�I:#��5��p��ID\NH�܌�-P.�k(I���;����1;8����<��Y�p����|�m�B��,^��4�Kg�CC�;F�|�������08/��mne������m��P��XY�	,�f��df&�C˵E�y��>�%�e��M/�	a��4���8Ո6��!{�Z��0��q�����GD�Wμ���)����j�~���~���bԉ��s
&�!]K��owX	M�'
|�YrbGG����4-,��+6!��g��rW��S�j2 �����%_O��K>��7�ʠ���Q^�x�4�� �6!ߠ��99��g�X�\La�T�%ظ�a�o��8t��W
ʑz�����d-:�@�澽�B"˝����e��Ƴ��U�C���D��TY
�Y\*�����3��4Қ�	�u�#/S/�Ѭ�"��F�IPL1ui*�d������T@,�p�Y����`�L����i����#�ټ��%e�a ����8��ٯ�Y�\e���=��N@9w=B����10k���3�"6ы�Yk)菡��|P�����Mz`1�aH��51"i*�e��7 +�s������)pM�t�(^��������d�2��@!d���� +�4h~�9�����7-ǃ?݌�T.[�XY"�g��>�yF@��o��`6�đ��G�}��R��d�xu���`���i�ub 'ljb2*D?wu1&�8�}��F��%#�:�
`��^�ko�d�W����L�)�V/��V�D1�\ (eX�7W���Wq,�Z4����5�"�PB�ry|�+��H��������
�|/�+uzt����1���[��k���;g1s��)!�B�cmm��J���;����ԯL��=O�;5!���C~�p-�nzi�������������9�����mCv8;Jy��]_+��Wϊb%���؎^�E�o�6��'EP��G��"i����q���o�EGn fD(��S"m�iNo�#W� ��}����ta�~4�O�OMvW!�w���.��D,�;��~�$a����̫��{����3�'�͜9�	d"�wܺ

d������u)���߅�C�I��'�a82sK��?}�'�(!S�_����,b`�KM�}�o�9��=�	�<BLEM0�CAt3��fӗb�zX����Az�W%�Fw"�oL�kj	�/�X� ������F�kW�:.���T 	�}B���9�!*�CSƖ�j1yH��!~	�,M~����3�L}׻����Eݦ9�V͇*o��8�@E�>�ׯŲ�7��j���ڄ�k����1�Ï�ub��^H�4"g���Z3$���m%P�L���U����4�}'�,�i�C�J���5���g`P(�4�&ڊ�'���vA)�����7a٭?¡��)����x��WXIC��.�ȓVC��]�5��U�>c����������7"Ik�@�ϛ˫�3<w��qՊz<��a�_�()���C��Ԃ���$\�}��P��?���rL���+�W.�Ǜ1nWb�=�0����[̿��'�DM�kI�YĞ��G�َq
�栜>����#Ƨ@��/�X(w /|؊�
f�S^
��9��#�+z�1���d����Ԋ6���)QOc�;�+���1��;���ޞ3���*#�k�H�AG��{�R��u�E�v�oOT{]0���D��^�����"l>8����
1�GN�/5A���E޴�LK�?�,���ٙ:dN�ύDi������&�$wc`��U)>J��B��^Q# �6�6��5��4�eaqu.:��o���?윂I+GN$����+&���<��ݎ]�1�_���L�B.�D5�v��*A�2�w��!ƒG�H�`�Ab��j�f*�:� ���.[�`:��t��n ���>�dJ�6�K._���q�?�"#�Man�aU܅%�_LL�104�J���Ct1�|�#b�3��D��x���?;",���!JV$����cQq/��J��=�E�a���� ��L�q�� ȃBN1x�I" O�w���Ţ*3x���]by�b�H?���@���r��a<���`P��G`�������X�B<����3��hǰ��
l=<H���e�"������;�E�M$�=y����q�{'���Uj���UF�Nq�W&0נ�Z3�g�&qiu�(���rj��r�aF��g�)C>:=�ݧ/���c�������MGj���E�������7�5<���Sw�r�,k��r�D�JC�l�x@�����. ��
*D����	vŎKg�����I��׋�$p7�MLL�47VTs1��)��V�����h����xK�{a`` ��'���/���&1�L��*��Qh����'�6�f5
u���$W�F�Q���i8=�'��|��e�;W���k�~��k_�a���O��� -��A�E���a������E3,w�������.V��x�¡ni����c��)�J�G����L�#X\����E5Z�L��B�9���K����Rּ`���Ԡ��T���n�9v��w�����N�˿S-��ݙ3g�5���)�b�͞=[���\�뚚�D�(�B�|nVx��? �r}q��"0E�m2mAZ����:��B�D|�NK1@�DE��Cl�V+@X��������?��.g�ěs���6��=�縮����s��Y,^L�6��-Vd$�u'l���ķD�e_�EK܌]�⫴�tOu����o�i����Z��������]�f����]�X�� q��w�+7(�j�R��6��{����������P���vu����E�Y����wZqM��8�:J^A���������0&+���I\7;#�b_��	�X� �{��>�z�~�.M����^�߃�,�7]Z��3��<�~�t!�q�J��u��!�� W1C4?O��B �g���$�=�nű��T):�T��[ԭ+��7��E��2��X�ĆJ�]�0�ǓǂJn���fƂKZ�HB�м�%y>��k0�"7��*J��i1�GŨ3�����8;]��r�T�g��Ti&fT�=�F�c��3HגˇŠM�Ϩ`�7O�l��̺?-��:�ڡ��,���w�=�a�|ihr��;xՅ��d/n�I��S���8Ol\�_l����	������WH&W7��Z�ǣk/)�A#	an��X��G�����Be�d���`2h�����zX ܨ7��0��3���Y �tr�����H���m�!�'x90g��@�K���ꪫ��w���?&����)��R|I�`ԫ0<��3�]Ƙ�HÓރ��M���'It�՚��7�8�j����?)��%:�����4ؽ�h����2Q�W8;({eM͚f]1ц��B��%�o�Bn��#S���1��$)�3����9.$Af�Y p���B�G <M�,�@��;�qK�	���=A�^!�I'Q^�
O0������6��W&���u�I�?�/��?�2�	����-�����Pd��N[.?O�'ujŻ'G�;>��<:��������L7MN��s��؈)6���g{Fq�g�Q5ZǮ>O;c����n ��T�
w@r�߃�,����
��77vG{ݓV���m�}3�t>���|��E%;����|v�\�ae�Gd�<����߹��e�;Ш����v����w!
���2ds"�w��U��h4�]�,�AJ����.��\��x�oi�*0�4;Cpgֈ�A;<�s[�t:��Oa�#C)}�~~.��\8� �d�H��fJ�U�j�:�V�"i�
v�A@M�rV��310>��M��N"��}�Z��㏧��qLaZ�A>ɺ��n��СC����/�In`��������=�PJH|������>+�2�2u�_~vM�^�����M�I�'���	OB����I�E�`�����{p.3#߈�h|C�x�͇�4��u����,��OG%�t�^xb�>�D��.�.D��?˘O}؇rY�<�y��h�y��������6�B�����)��Ţ�ab-U��9s�@����c��3 �9�`��F���͛7����𹭭��\E"�(++���?��%r57��!0��|�?�2;^��kPQ��o��6�P���'y�<v�5�i�6���6wD�@��bԫ2�z'��7{&.ǰ�x~+Y�aېC�![���s��a�Gm	�T�vb��Y���<��0�r�%yN��&���Nʝ�Fy.���yByy�ؘ���-��o|#���m�X�,�dl��W^y��7�~���rޣRTT���~:���,��۷�>gww��ǔ�x�l�:�������ؠ�0����8q�(�����4�[[i�|�/�������/�\���ф��®�Ax�5�[���+�'��?�8K�:���dͅA�0,I��KYbc�";�6F~v�X�QPǶ�����8k���늛)yR@�J�;��Z)�ׂ����A7ɔ�kqR�����=|����@��D��<8���D.�����g�K,D���y���L������75!޹��E����'9|��(*.��9��ȊE���ŏ��)��q�bL(��G,5�l%E�®kIM6�orh���v�J�);�nran�O�H��8�1.6�3������"-V����z�+ޱ��3J ����7)�1�܂�+����b��(aL;��s@f0��Ş?rG�K$|�$K���$#KY-=��A=%l^�{�ݸQԲ^=f���D˰O�,��<��ݰ��_��}���%�:��k���?�>a$a�q;v'o#��`��%�����~�áV��~�79pkN%|~q�D�]'�9��$eӓ;ZŠ�t
,�2��7����?�Y���c���©>	y�
�/���~�l#ӿ��kp�w�ũ�y�`���c��`Wd�#OG�3�E9�ĉ��$Q� ��`2JZN��#��� 'K,,<���KX6�ρ}��E+,	�7���w%r�v_�T��1�r�3D�UH$����M��=x����3�>�<�}g'V�XN���a��#��	���������^0�����:9�n��'/��"�&�Nn_Y�bA�-C#������z�
oS���mV1�	wr;��h٘���CqWǉ��D�τ��
]&e�!Q|�A؜>�R�	E�K�N��S5dA����,��������� �[��M�6aǎH�c�w���쿹��L��[o,�� +��p��J�:X�,��m�݆���ȕ�����'�r2@���=ѨLt��&lB!�J���cb�P��:g��&O	��炰}�y��ܸ�\Px�o���㯞�KAym��wBq��t����4�����<���#Ҭ�y�p�B�1{���s��eӀ'�]�*����ՂOs��9�F#��S��0��+�*e�[t�*��صkn���J��o���`Z�_~�8���ڵkEޑ��7�½�ޛ�i�ݻw�{O?�]!~�W��U����cZR��٥�h걡�4��"�8&,l=����(+/<�b�PX|�ꚪ��C:?��|A)�ca*�-'f��&B0a�2 Y�JL�|����Vʝ� ���^.73�Gۭ�ʊ
��\���'�d���+f���;0I	S��5���6[���t�ZFqm��ܗ�yoG*�嘛,Q3h��̚.<���c�&� ���^{�S�M}��T�%�θ��Y�g3`�s�5����N|Ŭ-��5b1'K�)�[��[��~��3$�x�z��lv�[Ըea���-N�1��ely�_hFسX��~�p�������{bˁ�}_ZP}�m�ό�@�&���cŉǷ�o��&n��&|���H�S�Ɠ���Kf橡��������!����bQ��y����(����t�bǅ/ę���ڹɍ��v$�N�Gc�8�������Z\_��Ms���BfN/��%��c'�y�w����I�:JV�%^���������67��O�+'w{������[X�Ȭ����$޹��g�,$� y�H?���-�z�����w����Y�ܘ5�߸�2셾�����ՠe�p��^��R#��^c�N��V����q]��7��^;B?�!ja��;e��h/Z�'E��-�፠o2gL�)�3�E.P��jc�`���r�6@�1H�'JVe	&��0�?�r�����#�uӁ��⭤,�E��.��}�x��P�N-ULo/[8o���f]�����Y�^�kGG�0X��T@xs]��3
��-��!�>?=��V��Ma�3x@QKQ%�,�B0���C��']��LBŻ�2�zg��V?lubo�K�a�Q�o�Js	~��0��#�sR�g!⎢���P�0%b�؉E���w0�� ������ҵ��
#}oZ�    IEND�B`�PK   .{�X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   .{�XN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   .{�X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   .{�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   .{�X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   .{�X+L$��� �� /   images/aad47697-5cf4-402f-a095-abba84463b41.png�wT�i�6��;�#��*��2c��T	ő�z/�k:"U 0��@�ޤ
��z���K�S���~�)���Y�k\�<�������~��B���_X~��������TTJ��~?wx�����/���T����[����j:QQq|���{�����,�tV�3sF:�R��h�W�VNƆ��|v���dq*�_�����*&a�ۙ3�%>�Or���������~�����~�����~���������~�ȾP��~�����~�����~�����~�����ʾ�?��?|�p~̘�����\���*�Ηsp��"��'�&�m��׳���C�d��;'�G�=�Z�(���/l���d
ʜ������K�Ͻo<�J0����̚��#�s>q@�}�OJY�n������dR5�/�|�(��'�����ȏ�c�X?֏�c�X?��k�'����?����=��$K���8b�+Y���L�ug��J$L�R�(���2R�]�������²��7�btU�謫4�
.=>��~ӹjWS7�����y��|K�]U����Aw<)�~���w���WK����b��yf_1<��i��\b��}`�/.o�U���(��ͬME�������Ͼ ��+8M���R���XP���m��FC�����Ж�D%�w��2K��e��7qoޫǉe�QfH>_'V�%�oכ�)�p{��ڡ`FS��GՕ�ᾰi�)A��+O�`�+�ع����U�&��:��#�S\-9l60�f}u�����P_I�?A��4�O�����#�W;:Hj����Deg٧���S9�C;�IjE"w��)���0	*0�du�K9>�~�\&�A��L�#��|���+�R},����qM���딴��e=W���a���W]zx��K��G���ޑ��:��=,��j*0���{t<H#f"��rT���
t�՚^'��k<�	7��xn��_����8´vsa�r� �߬:ۛd7Wmv��V�#�u/B橉��x�p��&�r��ix���v��Ǹ�#GY\��US����d�8�Gf�`S�����y×3���O
��:
�F��[��{�̱�Q��.Tb.�d��gh���Q��aQ�]��_��|�Ȕ�[�H{�ȱdo�7cγ�5=g:Ԕ�X�e�+�e��ӗ��ĕ������h
y�E�6�G�g���K.s@�'�K��Wk#�\�ʑ�5~�7�/�ݮ���*��Xֶ�1��\����xޤݮ\}3-���\�����x��~޵$��"y���^���=�}M�4�P���=H>�`o��9�/�k��i���#�B#(���z�~⍄��Edt���'as�
A�X�G��ZM;������{�?]�����	��,�N|9жo�ޑӲ�[��n���x.AO�B:�F��C��7�D���;��2+w�}����g��+��fHVotìkP���Â��%��a2�p��M�[��w����#�������!v���,�$�.��� _�����Y��� 0��uW���R�(RN\�M9� �ò�eūع�����7ޫ|w��v"l���ðw����Z���o�yb֏L��ߍ1Tҽ%�O����Z�:�*��\�)2�w����eb�x%��T�O����&γ���hL�l��Ói?�8�S�S�E�C������{p��s���RS������@3��9�j�㉪��5��5�#Q��gGM�\ݘ�v����;��3k�H�>��ZU*z�[�|��>ʾ�Ԏ�N��e{U��`,d�愈���(���P�lA��K�y�
N�#��x6��+��hQ�J���8׆-/���c�=�?4ݯ�2O�1����lP���[^�K��C�h�Wp,�*A��K�d�mx�N��v/�k�cg*��j�_��t�撃�	P��1��Ć��m�d4u��e�1E���?����~%b��m�����P����,�N�N+$�� N0�1�U�8�lX��vq#����`o���nkJ3k���A��T�L�<ذP��#�[��'�g� ��ڢ��$�ԕ�f�iZ�|?L)w�u����2�*�$t]e������"ߑF�!�g!)	l�kʶ)!C�C�jQgm�g�J�'��&�����q(f
v��d�H�^O���f��yL�����HeQ9� fC�Ͽ�]��n�l��̶l�Z�_�Ex�۽���u�)+�
�7��ǵ&jF���"*İ�Q=��"^����°1����g�8M�j��|����g3��>�J(�՜c�T��kt?O�uU�����Z�C��:\v�S=���	."@r���ӂrT�O���3� 2���!��y����3Uحɀ*]Hyd��/�x�����0kBɽ�9�)�\�5�KFM�1).f�V�y�+�[��WnV�9٥_�V��+ڙ�-�o&�gM��{�����!������z��X�Y��ײg2#�T�e&�:;���f�k���uQ�S�
_�j���パ9F�cL�Q��X| a�ev���_T{�+m=>d�_t�?���b�./$݄���S������8���O�F���t#�F������vQb�򕸓���=[�i4��û&���ڽ��,ӽ�!q�}��(F*ka���?dӯTu�5q`vZ���mp#�N��9��-X�*�����0}�������ai��Lr ���mWg���IYm���Z�=mRyϘ�R�4��A�J@ ��^E�Sl���x97��Vƅ��F�������zեh�I	�vt�P�'�%�lk;�~��ɨ���`WԾs����i�^N�ڍq�S^��x�O�)�%���rH��\���l�۾s���^c��OT��z"���}��+*#�K���-�E�p�5�j���5�+�m G�~q�G������k"��s�뙺��&.��-�ʷ���b4�����Gl`9�x,X�#,%������T��Y���<�e�ۓ�WR��Y��V��G]���eȗ��L��̈:��¹�fqoCMa��p�����-l���W� ��	Ѩx}Kn�JL����,����9�k[��z3U	-�w�l,�$	Ի熸 0�Z�	�06�G�i�s��+�S&���6��n��(��@��j�Ż��w��V����6�>q2���O��+��T&�%�n_ߗG���$�$B$%9��H|ЮEP�>�ZF����k��e��}jx`mU~�j�y��/eAf�)T��ؘ��ƻ�,t�������*aBn6��X��n��;�b���ų��u7�K
��Hv��S����T��	�t����⧖��
��,T�܈�ւ_�b�'��k�|���(�i�iO��a�쫊)v�|���ηzV�
�A��h��K�C�wQ�s)���(�+�s�� �2��1��{�f�-�}�I�"��`��]\N�co�W�������`��4A�z�T<�<5�u+�[�m�Wo��.70)Wǐ9w���5wѡ����\�>�6��L?�:'�|�h�PP��d���m٥.�GY�g	K��_��v]	�C�b��`�V����%/��O�灐0��6��O��9��&@��a��� 5��8�+��\�����;u!�p�P����H�i1���x����FZ��ϣr��H�J!:O�����z���`3ğC;<`��ye+�^b�!e�bq��O�t@�*L?�%E�}����|���ia�P��O{>m$�E�D?��ǚK�ӛ����$��Y,D^�K.A���K�[����:b
�B
pAׁR��� ����i�(@��7��z|���:/WG��s����&��CH�~�'M�;Aƍ8�uo���0����"����Y�H��^G�n�fN����#� �ˑf�>���2�c��$�54�����у��b<[$2�{�A�t��:��4a.�k:��p���b�ݖ{[�ࠚ�p�q$AN�fh�j���F.oA�rF�g������ �9�P��>O"��9^�Ɓ��
�%ȩ�#-�M����W'	i�\A�Y��$���΅*�t�"�E�A7�FRC�Lp�Ǚ9�+1�ϧ�����<�o?�Q5�����e/�pm,�oz+�ٳ7܉ÿ9k�E���s���Uɡ�!o�����]w!�(f�cH�����Â��a�x"�i%���PZ�I~��sj�N��7t��Q�X���������'}��ފ=�+@��=k��M1܌��u���Z� �_�=ߍ�*�{vR�v�rMF�)fҿ�,`�m�,�i �(| ����}|q�s���BML�GR7��:/7�^�d��I�:f���g<�,�-���.yC(��qV~�T�&�΢�7A\��Y�
��uQ��t��L/q�|�ZuR��WZ����Q��L�7����#Ō�e뼕�m*����w�2�)
!PU�/W�p�ȸ�B.*��ʆ�6��k������*3�O��B���tx����!�U��z�eє�L�c��)��<���#O|�h(��n���9hâ�ⱒ2s�����O��6]�A|����c-N\/��h��:M&�d�vg��=�f���}5�W��rf�Hg�IW�]�0Iyu�J�[���*����A2�=��,)�v[:{�i*�K���{X'�����n4�n�v����!YS�`�~,��aS���;�"_�M�o�I���8<~n�G��%K�7H_I���KT�v>iwL����r�@����6��J oĥ�|�Jz.14}�1�&�X_������WΘ�|-� `��az�\vޠ�u#MϏ�7?y��h󛼚oREٓ���W���v�>�boxSq�2�?oN앁��o�۰k��Cɬ�I؎�����^ �5WT�M�|��;��G���?�6"�B���J�wt�������#��r����MO;������v�n[�Ȫ�+*�9|�j�e%)mƶ�/|O�q ��>��W��')�z1�_���f����y��B��ч��4ss�\� �30�y�qW7�_��/���{)�.P1��0{����m���M|���y�uMI���zۚ�H�R��$�4Th���O�i�������/{ގ4�] �xw6�ރHʼe�QF�F/Y�ߟ��Hk�ڱ=�|��==���8�S���W����T��p�#ө~���]��aq�|�{|��W��-����!3�Iv���N���o\YlC�Z򹛗��CB�佅�YXގ�X"��ӥ��C~�9
�ט�L6����{g�����JY~*1zԜu�D�t�'Ɛ3ތmF!��$�莶k��N)~�� jM��J�,�l��h>(И7ׁɯ��+!˷̵�%b*ˉ�Y�A-�\z��@OO�F�Nm-�XH��VЈ��3F�O�*����"L��g��c�c^0�5)�u��_�$emo���,G�1�C�q��1�������ݜ�߈�(��M�� x�qlb�_m�&�w�5z�,��C�&�{�6*r�RU�d�ɗ��A�K�C���>"����_���ʯ��C[EY�1�ַ7�vy����(�;e�C;]�Z'
��{�ϛ�W�-6$C2�3�x����93vF�x�OхS��wk�k@8��l(��ǵ"q�c(;��S?L�6m,���0�N]Q���-={ �?l͠�6/gw�4g�+�F�<��μ�K��%%w���TC�n[�|�������ea?��t}=E�-��_z]���kf�\M~h<B0��L�HL*�o�O��0p��.���f��EY�&��������oQJ���,���3d��'7^IA�XoCO�#_Y.�S�q��{tn��2?���p~�0�����w?gػ����Օ]��`��zKd�d��Y��r��#��D�h$��B���=���Kx	kB�)"1�Vy7=g��z
Q��V�=?=�LHh�_r���"����4�B�z��U��"+B�a��o�Y���>��c������ʅ��=��`�P2s0�q��av�z6��m����N	��R��E��a:#n�|9���\����d�'��Y�\u;C-�A��}��4�X�r^3�S�`ʐ���Z�Q<��5>Sb��X�EH�	���~a�DW/�d��-�ŋ�$�ҧ�i9�k)�=Վj;�>麨�1�Д6W �x#r��s5�3u�B��:��w?}���(Kj:�
���U�;~*Q�t����B�����b� �mx�	t���g�m�r��r~8�`��cJJ)7O������V��͇"�3���^f,�>µ��H���O��H�B�Y�1���x�O�0�)�:����(yM�s�.)$�ZC�Ȭ����!��Yܧ�3v���s�7>IA�p+��nJ�`���p��96N*��Q/0�j
�ǐ�fZ1��&��n���W�{�ǲ3���1Z����"�k�!�>C�<�K�Wz�7Nv���«�tbɤ/�")�aw���D�鍊g�,��*�IR��_���Pl����^�w�o*h�x�����A7N|~G/����o�f+݁>�R�d�d�-��d��R�OI�ba"��]&M�o�����OJ�ӡ��[&ꊈ�Sn�ʦ�d�����qrJ�I��K������w�f6�TE�AG��bPH�<<:V.ܺE�hk��cM9���|���~�XS1�C�R�2��^3�}����f�GU��cц|��Y(��+@ 	��4n���r!>���g7��|%8�ش���1����4��TkIg;�c�Xw�3ۄ!k�-��lo���C��0EE���{�!��Q�������cI���񳧗�tVlI�w`?�ƈh/���H�m-qQa�ѵ��wBt��. �v~����������1F��]_��'���E���ψ?�'9���J��,Z[��Y;+N��S�%�����[tE(:8m������g�"�hE%s���z9AO��۵R�֗�/� vW�O�N��P9ϝ���Ϝ�.�Ij��,oT5����bo\v�`�)vk�|�9��-�||_���8������ڊZzyh�G�̀��=�aŨ' CJ����E�N5ȗ�r5��NN��H�.��5rP�r�Bȱ�
�c�R��O��|g9�����BMTH�P>\��p�ˤ�@S���NTO�$�R\ʑ�.��8麆E�e��1�����d�� VyƓz�i2��Iڐ��a�ZJ)��P� �%g�Zݶ��A�gG�w�h.hc��L�~�˒�_������^y�r����)z��U��=~����V#���Az>%���ҷ�(�&��(�������w�Ps�J�c{�G	�5�F�v,���kP�St*�m��rJ'[��Rm��������h��G?�Ÿ��ny��n�H��fr9xG����
���}I��o�*=�F�[ ��L���|z�"��E��d_S��!�|S����'���ә ����k�����A��-�:�Hs5w�IW6sY��H����堯'T�"�"�6�7<��I�zI[Hs�-n5!��+���Ch{{˨��;y��$�.�5w��M�#/��3g�2�[����'�R�y(mSe1���}��x 3^�X'
T��[|�k�Y��IiI��ꊒWO=������6�{c�xE�p(��Y��J-#r[�ɴ�������)�3�.�sװ����؄�ն�N8O����nο��B�� �d@�+at�qeȩm��B�^$�Ԇ�(��Wi;­":ʯ�	��i�(O6l���L���6�w�P��l��V�w���Pf)���D����QΫ*;��#݋~��.-ʹQtvl�,":����{T�� �0��d�k:���o�`L!0��0���D$����ֺ-4�44�jܫ�M0?�{;�yq���}���{,�ջK�c�[��[���]g���OlSG�Dj��Mh����+�����f��
J�?�'d�<o��w���}��3�*�&��j
��g�bsb
봚�q��kO�O|*У&G�J�+����`Gw�j����Ɔ��>�Ҋn�<�����c�ׅ���;-ꗺ�%�!z��`|.9��Վ�bҸ���̟� �3�t�EڕECA柡�1����9!�r�DOM�.���"(�n�JTey8Z
���˩�c6[�ō+e=����FĦ9�����e뱱���ǯ��Y`�Hx��9~��(K҆��`⪥��0�R�N{k�L��wM5���W�Ym������G�Wd�|�o^���M���RXH�%��՝B�����!���w_�mnV'���f�� w��W�ǵ���7���cY��r-�wJf�h�0�c����I*���΅Z*�m�H����'�ls4�Tv��P0,�'ꉢ���`���w�`�0�;i�+_M5��2�2�{�x?���/��|�L�e[n�@8u�.d��'��4���h;����F{��8�%�Ks+1��Q겨�6���O�[��Qo	�l��� �B�+�W�xK�I�u��a�R��7x7�V4ὣ�����/���Sni�cG:|�\K�����W_WK�?R���([�],l�3rMĊ�ڹ�юV�]~�7�@C����?)�`7��}�T���}�,�#$�$Г����N�߳���e��=7��|hx���w����-�"���T���۽�Ǭ�F�a���8�Kz^f���irճ�(��_f���,U[�R�`C�E@C�qY�����ShƸ!�ɸ����_8m�aF�+��a�]�y;�a���?k�H�nh��aޓ:4�	��oIc������� @6�oT�Ӥ
�;��a��p���9F��cu�y1HQ�٧o%C��@q��Zc���3N���,ݥ�Nq�ec� �ym�Lڥ�j	r�A_9Xr���b㸫�0�Y 3I�������rJ�m^J77��m#p�FRB�������3箿�녲���Į���B[x��~ ��P+���-2v�,��@��]�ud;�ٰ���X�i�����k|%_��|�L0�E�jmNv��)x��G-��m_J��t�*�ɻw@~�q7k�4k�iԕ}�l��43#�����aJ�z�צ��~�;RmI.�<9�9 ���pȉ���8���h;K�t�I�z����fRT���U�c/�sM7)�����?���ƹ��N���L�����+��H!�dm�����`��[2 $��U�M�D*2ŝ3)���n�=��xu��pΏo+����2$���eh�z��`�J�ӚL�>#������;�����J����N�S��|��-��'�F��p%�&K���#�3��)ғա]�)�׸�O�z\��F��D�.ϻ.@�QDqe���؇�������؃&��ͣA��k7W����Zqc�����5|��Z�gQ�C�"���������,=Y(���4'��JD2ڹ�{Gpeʕ���.T�x��e��q9���=Ѹ�� ��`It^j�U|����6 ���8����*�`���}���3�R�I�X��/�'�zH�phC[R���0�KPV&Y7�"���ֱˏ�% ���r�'��\��T�^�r�=Ĭ�3�U�P���f�NT�؂����*��6j2L/�P̡!���)��Q4ԒzAT�T�wa������	����MF�k]�D "?��4�E{�a5�e�Ԡ-�ܩ@�R�u���ĄV���A(�^������&}�@���dN��PkY8fVa9������	���'	%��\YUS�Ͼ�eOW.��2��^��B`Dw��t�wA]�{!\�K�}N���J�tN�ƶ9�4�)B8xB�dfo��C��(3�/�}}����'_ٓ&i���|������^&HzL���pB��Cd�D�Y���3����=q�;o�U�������S_ QP�{��:雏YuF�����5u�������NO|Lg?5֪h�V�67�6�p�7vPt\ך��=3�@�. W�%���؂*m�E��Λ�*���P
ʪP���`�
�
�qN�e�פ�<c�#�y4or���Gib�IZ\��[�X�-�Ĳ��,���������o�h8!��l}��)kzZ-��9��khk���O�	PA�\hC��1���3V�>1�����������w�kN��#�Fi��t�S9������/O(�jm��3o�x����=�v��QT|��϶?!m�2��IO~E�	�5ƛ��`�7�w�Y�g��i%2p8�Z��nsp��_<�fhB�VR�=�e�S�[��?�4����5�B�ݎ�'j�{��Z��x� ��'���2ɯ�N�2�g���]Π��`�q>#�Dg�,w�j�r�Hh�o�FG�ǟА�
��s�^��p`�J�:7��,�MT�r�M�e��Mg�~b�Z��}�Ŋ���4�����*e	����ӳ�5%������I�]g~�O���&�nڦ��c$Ռh���/�MX�}���s����U�=K�ܓ׌灋˂Y���c5�m�&RP3�t>�.�6$��Rh�m�c��w��4�d_#��A�	���[c���'z�ճY�f�pׅ��,�GP���Du�DGO�g���:��2�\���0n��_#ra�J-V����.��{��Ql����LAV牓G	I	>|96L�@V	q�;ܪK�m�42���L(xV(��Yr��m��� lQ&"Gʶ;
��?��@)��5�Y��me��lG��~z�{�G�F2U�n��A����Pd�k xkd��(Б��tx���]��~�>�����q���+.<y��fyl`,/��{�a��f~\�]��+j�����KO��͎3{�if�W_��~��/�3X�[{{b;(���<�G�uj��L|&:<Y9$��Iln^a���@,�ns5�����?�'���LG����^��Z-���\ʖ6Gl���N[���sT>���m�C�f��j�3k����x�+!ʷ��Y ���J:��r�0Fذ2�U%���/2i��::�R�=d��C�.s����hX�.����������oΜbH�]�P"�3�OOS�"�8��o#=.;],r��@�!Ƣ�H�UH�����Z��B�4���^��:���3X!�Yx��`��Hi+k=�r��)�dA%�oL,Y���w��@]�zڼ$�2e�1j0�����x�jG"��ڠ�\j�m�av���D�fGG<��_[���Q���Z̐65��¬Hu���2_�[p�T�S�7�3-��I�w�y5�o��y������@�5���y��*ooJ��U�Ie���"A<E�o�F=@]�'��o) �,�㙜p����Q;��t�X!H��ǉ�����\ȫ8��4��=U��<9ꈫ�+a�C��b�Ni�%��#��Ѱ�2�H�k� '~�k-Vu<*��*5`}M	*�8>~/�R�LG�R)�"���u5�͏���F>�����A����!�ȗ��G�0�H�.xH|��Tg�[�6��b�.Z/�uZ:@z~�S�����tE�/����AM"�au<,�wH�~��
#���CǈybQM��!Es�ᶖ0�3����U4��$U�������{��� ��C����M7 ��X,�K�nS�܄+� a��!���ƚ���,60M���w_���_��Y��cz=��~%)nx�Dա�l��n=Dt#o��q#� i�G��-�y	�T���G;����2�U4A��ШW�'�>yr�k��f�NҨ�O���s[M�������m�g��Dq�҄Տ�q��7�_G�ԃD��5d�A5�t���r��`.S�]Ͽ�S>PR�j�u����\���ۦ����5'����d�[KY&m�]GK#hZ!�[�s�g�jX�.�������������b�.{��=�!�> W��1�8�@��R�j�h%YY��2,f�C��C��՝-� D��m8k����t���>�0�;�TL�b���s��Փ-�7�&����r4+�y!3B{��M��%�駠}�ųGw��".��f[6/q�3!v�DW�+�����m�.�UA�?􎅽�dn����V|��)#�J0`&|���A��]ɚ��ظ�廳X��&E�%:�������	��ꏧniIp�D4���}]/�~}�5�3���,�ƾ�د�V���h5�,�Y�۫�f�^�,g���g�	z4'kT&�/]8~���u��O�k_
,���S1+���O�{����yC��8�xt��T��xV�	��5d�f+� �1�F�W���pD��q�N� ����́)��+�i/`�B����E�:����D���[j5����g��3@r�'��o��I�t57�.�ÎDeFY���uG/�zrC@{�da+x��=Լ��E:��/�X��w�Yɑe~x��K�b�ʥ�����*���ɣ~m���88��7�Y#��P�0��BF��^��8�~������M\lP%��W�@-<G|���̾���jw�E�w���+��Y��_�{�{q���ˎ��l{?��=Vj��2������-���z�]���%��n�����z�JJ���ᜎ�����D���gB�Om�f��s-��]=-����K�Y��h���Or��Ǝ�Z,2fJ�O�]�����Xbи�d�׎6���J�,{���}ח�Ŀ<M�8̘,V\��,�݀�ߞMY�\-�ag�'�{%ӳV��5���rbQU��j���i��MX�o��F�M�!��\m4I%����#c��H���z+����k�C�Pvi��~@�N,[	.9�U�1A��Bw��f���|M4*��3nc3��>��3����Ab���Ӡ�[F�t�������E��B�@tq�Sj��8x��DRDBD9����x�\�!��� �W��m�g�¨�~ٙ��:UH�~�n�|���$�>�U]� 8Ưd�l��)�Oו�JE��⪌��������C� ,�hD18ΐ��j�"����c���`v��J����ma˚�]R�������P>~�q{?/�7���r��vi���-�����&;[ړ�L���{��cu���ǌC�`p'a?�����g�������;�Ͽ��Re髷l�4Nو�X��,-����jl��=��0l����D�(7^��w6�I����{�%z��J�*�V��OɈ�/�wrX�^VƮ=��o�^ך/�L�r�S��B)���)*y��W�q$�l/�}&{�[@����z�%V��U#�6�hm�簅W [u�c�G��\N��_r���kz��2<dw�*�e'�q�%k�/9�b���������`���Ÿj�ib����m�����rS���'Pg �˨���xr9�u�v3_W���� ��bA�K��2>v9�H��5c���?�QG�ԫ����v�#�F)�kV󭔸>���M*��*�z��.���>G�t_�*ky�u���H�T��<�1GB^��H�y���}��Q����[v5׉;�`%x�ؙ<m���v3'�7Y�����_�e�m{��6(]�fJP�捊�iR:*�t��g�s�g{N@����5���&)K|a�'�M��HE���d�}�Ez��\��1����c��j�]S��!������>�1f@�%%����z��;��`zz�z�lQcM̛^�w\��D���~�l�8�o%�@0�n�Y_�6n>��mhD�t�z�.l�$ �`(.{%��)U�t)mF2��o���Ãs_���Y�Ð��Yw��3J䪂���ցd���Wm����׏��\�#Ս�h������s9��ݮ����ݴ�,�4�P_�C����m����!{�	��z@��:�+%�K1�RL�3T<�䷞��y'��u�p�8Ǉ&�^��O�O��xiu�1~h8f[�����3H��c �M�W��K?.���Zj��D���L�z��gd��q���y�h�j�qJÀTe!�|�����i�
Rf�N�t
1nPS���nfꀷ�r�8�G����h'���e�)}6�W$j}	��[ �Ç5wP��8���㜕<�w�詠k��,���7�=��y�����*
����l��c�� /�
�M96U�k.b��`�dQ=���)V�5�gUl<��^�F���=Za)�n�+)͔�h?F��<T�2 �!Fo@rw���4
�3��C�`��ƨ�?ap�zΜ�k�jljѳL�yx���v�Pf�����N�H� ��/֥i�������ԏAId5~�$���2j����C,b���;��>�?�����q2�������<�pqo
�X���Ɋ�#��*P��6�S�, W5u�(Ιl3�=��5�wc
w��L��V'���QQ)��hK>��֮ >�w��Mwn�
�3@�����q��q�*]9������4�k�{�O-�y/�G�+:�Y�ZD(=�a��i�'pmk�P���bB�6k�J\Bt��k�oGx�^=6!�G`dEĜ�E���-������\H��������8�N���h%���N��t��"�>�9�Ɖ9Ip��zp#f������3��n��&¯�P�!��$P�����x?�����ޠ�5���Π����������?�u�לc6f e*����儇_v��ٸP�YK˕���GgRW�w5l�>��·�M|��l��(М��e%yO����]\BY.�]�z���7Sc��ٓ'�f�:}�jw׮_�J���-om#5i�*Ė�N�>L��t��>D�9jY�R���bjzM��㷵'���=����L���g��V��H%����O�:Х��>�F/����Pk�f�
�^=!�)�w���Q/7w]_Ջ��}_�tD~o�6��e�bSb�OSNo��O����zj����Ē�e��M|��j'ܓ��5�E="�T5ʞ������=�Jr�Y�;����[���I��9���C �mi�T>�Si�y}�/�R& g�Z-}%[~F����m~�b��|B˷m+��4�*�\�q��+O2DA���ة&h0u6NR�{��+,��s�=�/J�[�t�F����=�ua�9`�l!Ro��y����݈X��f�5x���{p����&��RlA��F�c�#�\��
�|<Zʥ�}��ҹXn����7���_7Ou�a�6#al�d^��(���8/���ҵ	�5�Έ��8���5�L��;̦�Q����o���V����1JzL�zx�&0�ť�6�aa���C�#��<\��jG���^)h��}>*�����
��m���R����'(��g���2R�Zm��t��[��ֿ��Al����o�m��5�Ey���]��MC���� 5��G��u��N�����-Zݭ�v,�sA@ y��	��0I^O��g�vx�O{��p�s�pjM���A�
��1�G���ذ�_ٴl�C]�{qGF�(ag�
����8yt�|�'��[<$h��>����&}�sF�6��]����F9 ���7"�[j�w���U�E�_<�W��
K62�lɣ�@�w,�z[97 �������?i^�hBHKL��BD��N�s]�]�;�wR{��8+F�@h)M�-�\��4�-��v%�Z�Ҩ'zid�o_�83?D5���&����n����N�%Q�e��۔��@H+�C9ȫ
|���͒�U��Z)�3΃1�'>�f9�Wtf�Tz	$m�q��LZ�C<NF	g���h�&�sR�z<�$�s�4-�)���:Z�u����}�`����曒ݯH�k������Djl/���yos`Llw��#��R�Kѵ�Ո>�'�q��s` &�o����r�i�0@��*���s.
2_�%��n��O֭VVR�F�!Iy@�"�m�kjV,6S�G���P��j'R�� ht��U���ΞϏ��sn�H*%����A?zt��l �ރ�kv$%)���@H���LW.~�YV��iп� �5e	���8�>#�G�6sdX/����\[n�O_iS��#B���0��̀F~+��̭�|�u���A��/5ã��w�A%|�*�9���O���?�(f�Y��X��v�:Y��_�E��WO�]�������*2���z�`������ snN�M#;��(J<K��pDS�s5��ZW��<	WtJfW&sL�p,���sOree�D�h�}�:2����FE�W�ֹ2z���n�^B�3Z喖=�je��#�	�nΘڠ���UFS��J��ѻw��<-��͝�J$ �MzK��P�x@q��j��|�1�ܬ�'Vy)(^��=z������10�M#�c�i9m���J��-T�>��/t��t�=]����gD��,�򧙮����|��c]�u���@��S�瞵5�]�����Hv`5��j��h�N�2�P�����)+(�o�}5�|�!fP�N�<�q�RR<�G+�8�n)��O�TYQv�4���A�$z}|��xlmE�[�Gf��/4;�l�ύ���N���ʻ*����Iz��:�7U�PUZ��s�œWfT����'�kO��X�t 6�̫��
=��ڝqx���� �2�Q��Ҹ���5ۙ�B��!�m<Wj*4��K�D@����}y\��
U�g�$i��G^Mva�1��t /�u�M�zM\ q��	�_��8L��ʏ�8�����<�{��7[���"����#˩$ �l�q
�����'ʋ,����LP�ʳ]k/�:E4�k�u�|���U��2�Uݨ�Lo8��˥��x �0&�<�P�Rt���mfU4�׳�g|LM~�I�*9h�� �fA"%@�����>����,>�ZP}�܍ O�톽���
�ɞ��w*�1.���8��W�׊���-� �����t��C}ׇ_Q!�O��+6ˎ���̀78�}�%�:{d�r��jRb�G 2�,�mR*tlxY��2�Dk�+����潂y3o~4����Ti5PLC��X%��x���HpL���K͖ ֊c�u��U8�[t�"p�z�֒��<�
��[��#%7��͎�����P���}=os<c���p;f�f�wN%~���c;���N9�̬I^�(�X�d�[��Zm����$5a=�����G��偁k��h�F��s���j+R���!���1�ׇ���3�T�ż�F�Y�Z��^�+@_S! p���H\u8��bN�Vb:f�T��jc���#��_�(�3� m<K�|?߸�pf�%��G���ʖm_U	�^=b�̭�]2�R�f^�����nD�]g�{ZTBl�ԏ�=���M�d�`o��(/��v��d����!�-�݂،0�����������2]Bu1.&Ք�ǖj+���=�^�OO�6�}�^�{X3��"3��s1\O@9�H����k�� =��L��d�[V��U-4e��.��{"a�U�!�RJ�PS�iT�G�K}L�$�dn�l��YE�/�A�-�Ԡ�ط�L��\����1�e�}$��'SK���'S�yjc������|�zm���S%w�D
��5k�̀#���ɠ�7�n�O��
UǳL=to9�*v�&��g|:�027��[��g;��/�_S/لz��m��b���4���_�)�@�M�V�����RL���I��!�=��	t�x�/�_��P���nM� q��y<�P�wW(60��mKm�k�0�sã�kFT>���.W��cSY���=EQ� x�I�r����e���R���5?��q`l��ȵ�n����q�JuX��T�S�w<"��τ�Z�~ex琊jO/��,"ȒLg`���6��@c�` �/'���t�ݹڶ?բQ�ë��P�ށT������T�]YY�ܥ�$١��E(���:�cӝQY���C�������{�c��^�����~V������z]
�7��K�k���@��.���H��۴�C��":ǎ����Q!�����jҬw�~��s ��ot�.�:�.��[j��7\��܎�p7L�����:�? 'R�x/R����Rݕ���[�>�1����C�
)�;L�R^���+�����=�I��lzw����s���-��2��K9�8Vվs�hT����z�����>�
�2u02�;��w�|�k/�����2o����#�/c�G�L�6�h�:�D���'1 ����%���)/��<_ � ��0�>._�Ɲz�O�F�\�^�1.(�fV�Ր��V�pؼ��lg7�b�O�'vY���ޫ���}H^_�aMу�K;s_{A~=�}������?�3�wK�(�h\R��	&�1&��=��g�]}P���]PVy�f�����E9���4�S�O%����٩e�_�&��̫ϵ(�0���*��?=�u��e���E>�$~+E��oA���yB �u�?

����go7�v�N���	Q��,�r}1 rt�y������ �;
9�%:��8�15�=�>�$��"��~Wp��}�ܝ���W�	g�	@���x�����S�.�w�z?Z���{�E�5��`���u�d��F�r�I��av|�^�y !� L��cL��]y��RV�b��h�o��Y�=&����2����MB+MC6ǟ�z�MxI:̴߿�v��`��{�<ψ���?���0��
��6[���?���)س#���9ɼ\W���pPoղ���o����&>P���qQ�D���n��z�3��-I��c�2/�ʞ���%���?k�ﵫ�[�W��×��nC�wfe�I����N_��,Q��QbY#6�"����s�Y���t`#���*�N�-�����(�`\":� ���-����g��@�I����Xd��mA>ݛ�C�� &`a�N��"�La0�k�JR�"e@3�z���8��������{ۥ����U����Y$���ֿV�e%y����M��`��s��c��M����bΝ�1c�8OӨ!�o��=�t9�+���o{� �rg���Qw�����c�
<��lvǝ�3��ƀ��_<z����F���9]�B�7��_݌7��Y�lɀ��}#F6uB^�p�ޡ��k,��M���c��CW�v��=���Eʖ���u\���з1���Ą�e�pb�Z�	Xjc�;,
n��Pޥ���VǅәvQ�yݢ0<Z�M�U�@/��v,��7B�a�d�F@r��{��Z�2��f���?H���I-����YxW��5�*r�⸉����Z��Ԥ����=@�����>L���i�U�8�s���j�FW�&}�]����� �I?�
&��'#o0���u��!�K&8����)�y
��~a+D1��c�ɕ&L�o�I�4�Y��?�uI2���pպ�������)���gg �����6�8=`A��%���j���8����Q��r��m*X��WS�6ʊ־��2�E�4��!�{���怟�#s�k�K�JRNJ�>��`o��|�w(�&�+�?ʓ�gTN~r�KP[
-W��6�rfT�g��"q�z�*/�k�'BW� �����5bfT������#�ɪ�Bo<�6Ad��%�fv��vl׮��P�$t�����냤���Ñ�N xs��D��^ό4�=܍$��m���m���mN7"\}9B������6�F���^�2Ň)��=�3�J�qs��L�ՈW�,�I	��rK����k�����Sr�6~��ki�K�aj�)� )�O���\�L��|�ps"�����n�����ZX���f
;��7HW^sx�;zb�i�+&=��3�=4%�����e3ҦO�۷�<w>2a�"z\��{P(��f�S�H��YԄ@�d��Oxt�C��%�I�f�~�JP��VLM���#<���4"/�R�z!}�!'A��)6Q'���s����YJ� ���:�ݫ�A�s��`�-l�#,jc��%��b�G���L�� z|���f-Wb��8�iO0�
S���4�?�R"���/��ʮـi��^-��>��MB�j���gApL$^{��?��ln�;�}���X���4����^��p�h�4f\�L���$Hp�~����騛��(�q�Bmǭ�z��Z���C���P�B�.��{���B����R��%���fO���']n��g�U��4�Z�p�5��N��/w��Up ��z&�U����nCyc(�$��g9W����G�{�������;࢝q6�'�3�n�ìAd�>=H)�:.ۏ}Ks
�N���qK�u�+�-�"��۩�_��'���6���6��Ƶ7��4X I�/_9���+��0+���ejql�hsd����l��ݍUwS*�ސOc�i�_��hg��1�~|�E���H�|,k��Ĺ��VBwK����FB<�f���jd���|!�a��-PZA���sa�D��"�SBHN�ﻙǍ��~��8��OcNri�J�A��)��*T �$46�j��U>cu�P_�l7��YQ#���BN@��en���+.�uE�BS�E�E��D��M��k�����ӯ�U\a u�+n��/,d
+8�i|3����\l�w;�{��*��GV%���+�.g�B���b�I�olnpE{�� eʝ�]���W�w����[����!����!�Ғ�'Ѷa�	�4��<+2di�&�7�X��+��{�տw�J����֭!{���E�R�L�����9������z�о��>D�[Z|�X-K�;r�Rϴ����0g�g����6���i`1h['��,�G-�2�e#^�ְ����[���aL^��[h��Z�?i
}�a��Xv��kz��
ĀV�%��#��G���%����.�g�Ɇ|����P���g���}��݀iL}u��m[�`��H�B�z���n��v���� ;S:���C/D�/JX,���2f��)��9~�k�:���.��0^��~�2⡤�T	yI����?�FE��M�r��D����uc���r1#rN5q�B|�C;���|��C��i7Z����c*6v�T��w��wyG�Z6SY��}�#p��s3��`�5i)���Tx�������%_�e������3���r��������c=��!���x��_��2��m���P6����U�K�H���^�r�hk-�d�}D�����bq��þ$F��Jk��75"<����n�)!2����o_���6W.�z�vyV���%(҅��[����-���:��L�V�b()a�$-���up��oE�F[�n�k\\|�{Z����,hi�vd�d 4�N�tݮ�����u�v�x~� �hI;�~�ԣ/=�m^��1V�&qPc[Ϋp�-{zSj5���K��{�}�)��f��Du�L�,��]���n�,���`��;3�GO����`��;5V�����ln'%V��h�_?��&rh�R��:�]�����'Y��v4oR!�vǨA��sBh*�ƞC���\�ʿL���hp�^����)H����U�� ��=�<&M�v�_����8|o�pX,+���҄����,�r�WP��Ev��R���-��0�5|*�{��:�=���`Ux -s�����P�a4�fxز�G�G��4�Qa����9��'���HP��{G4���}�H���^;4��������h�2�i �|�H^�Y��r'{RZ����ɜ���yx>u�VD�
 *YǳomA>A�	R��g����P��x��W-v�[l͋�͕�q|�:�9�?��?�-X�?U��C*�a��T��N�:9��M��f-�q�@��韈�81�m%��
�K�1�7��z�+w�G<�3"J8C3Y��@�U�؇?��Ѓ۔�P��Y�[�&7���Go�yZT��]%�g�?Xw�w�2234)'�ΝU� ��b����gC��o�ϼ��z�k4j�G���ĥ�:�����i�z~ކǺ=8$�,�@�N�����Fj�w��$~l�VG�Vp���*����ej,��^�e5�k����g��8ۯ�."í�	�k"���_`��W�a�l4����d���~�8��ʣ�&f.��>�����
�ވU'�Ӻ�R�r5n4-vhf��G�,�������ЄC��h/r����ݲx)V�X+ɭO��®�T��x�p�@l�����=F*E_w7CEK$�H;`�5���!)�K�U�}j�Ǻ9[���*[��6#��a۫�AJ��h um
��e���]�'I$��O�P���o��3��q���e �
+Wǘs�Q��߼1�L]ݑ9Ԙ�$���+���WC��2c���ͥ�]�.Jk�{���EBR��Q1vL���T5�ӆ�8����g��?�X�����������X���8�6D$��ɒjQi:+
���Y�KO�];��F�����}N�Զ�p�s��x�9Ah�w���w]NU�l\���)�*��?����Z�=������Ig�﫟	[���@su�CF�. 2�2�c�C�&���@���ծ�Tp]t��al�<�?mҘ0���A��]��<@Õ@�,�M�T�:wh���P���
(37{!��M����l�1����u*���T�o�xF�\��\��b�b78���R�Q���c����;K��Z=ɖ��$��e�Ԫ� 姺쭝y������g������!�jO�Zmb���sd�o��-c�q����K����'^��0�sI���G0xÏ?�2.w^��+���:�\�v�g�W-@�<X���,ÃÈ/ˈ;�Fai8��s��1�m�0�E%D_�b��C(@� 4�HK�+�3&4������B�* %٬�:�lJ�?��Q�����p���Ѫs8�ׯ��{����S)�=�]�̮�'�B�+-��?'-@���s����v]�Y��3B<�_�j6�g6�L=8�
d�t
B�Gޔ�S�-a�J�� ͒&vv����I��0.��Vo��]�D�82������!mg�����+�=��ly��T����B:��eKl�,�-+�K�Gc�^}�t(̈́k���M�q[gש�u([�Kv{����8&���s�y��< �(�1� V
���W�N�����g����H�%3� U�"`�g7,5Z�xlV��Ց��ͪB�
ڢ~ێ.{��50�Z�l�ŕ$>��Z8@5�,���&ٓ���sX���$�D��ō�H�C�nva1q�/z��O��y
�[Nu?�W�Es�ΰT�]V��o�_B?�6_�A�1v���J�h���ƿ��Q9R��:8ד�э�h t;��8�l��\����3��vl�Ƿ�	]����;A��D���q��s����dcݽm%ԐZ�gYN��k����#�=����|�ŵ�
���O_����ڟ�\���JI�����Θo�c��w�˕�*�#�}�����Th���r�O��-�@'%6�
&�K��o�pn_�f��:��?9�oc�����<v+8�E` ��^Zz�ȸRh�~�� Ԉ�������v�<� ,�GyG?K7	)�ѻ�O���uȶ��Ӕ�����U�0b���M��L�+�ƁA���kV;�J�g���ߧv�����E���~�&�	�PT��y�����h�з�fhg�C
	�[嵢�B&�g".j�QHo���A�{�ʹH�����
��ۥ� ��������+�UZ������0��,�&�ρ�aL��<�N��f�~�*����Y�M��W�b݅FE@zN��ތC7iNsK$�-֙�0�����jo'Pm��NBj.>������_SC�vP>��R���ǆN���Vj���7%��H�O:yW?��`�|�.����T{V�1�~�b~
��wa�0����9r���g���D��=�"�l�����\�����o��al��_q��fȯ9�F����I����o�PZ9���?wl�e��e(kw��v}��ؼ:gn%��iɨ���a����il��̧�o}�<�<�t_�(��A@������9�K����*/�����b9�<i;��;��'����i}�(l���̩v�և�J8`�Dfc�h�����ꏓn�UlJ��/'?��	�Q9�QU����~��S랠��z�|�-�p_n3�6&��a9S7���l���~����?�`cZ�`��o����>o����\���ѽ�����yCl�
(��ˢrq��}�������;���Zfɼ�]�:�`����²ژ�_��,�@�4�e�����a�uVH"&âfl���RN�{}��q��6���H��E���3>��C�'ݼ�6��cs�W�i��lZ����t�F����0��:8���;i[�;:�oµ�wٮ��3~|���]�ZW�K���!�r�,�	�Bګ�Ġ�^���Gu���V�E,��s����`c�����"���ؾR����r�r���`{H,{�z�����a��q��AۀN���Y��:��$8�&|�~����Nw�͓�gX�g�׮~ϴ_����|�g��R1�Q�	{���w�����e�@T���<���t�]t�����hu�d�8�A�I>'\ @�4s��W4�>��{�iK�ci�G��\���T�W�U9Fߥv��3_6@��~=h`���h��PuX+�����"�4^O�ߕFK�w�"�*)����Ӹ8�����\v��l��k�&�[B�����۹8:L��o@J0R���aƩ�l����83'��6 � ����	��,{&�Z�W��TY3j�.,<p'e�'� k���|���r��'��/M9��pɛ���,���A�&Q.�2����3�hg��j�m�I�V=���t�\��E:�M�%�n]�S�е�.=h�l�<&����\2���j}�p��?4��>���$��>�DVIs��o;{&��]�,kbZ�Ǹ�V�b�{���i�N�]�=�a?Cc�J�k{������֘̐Wj2]?�m��][��t(ЪĻ��E	�uNq�p���D�CY/@H��c����v`L��z���>��y,���+�^�dP�h����	ԓ׭@`�Rd���$��؈K���`�v1?�*�c�����[�{��� ��P)�zx�=]&�*�Ze�	��v8kJ�H��V���Y!��Clܛ���.g�;¨�eTo����,�=G:���XK�!®����s�U2�r�d�-�
f�a����<�3L�C� �Cc��>�бس,-���V�Z�������3	����{�jl:�D���VΫ�(�_
�85őc��r! :��k�I�5h��+;�H J}c���<�������8UhS�
Ģ*�U@D��y'�8s�c_�}�L~էn����Q���ߨ���z���^",�n>�To�B��ͲvJD��ݫ�% �o/�=T?�Ϡy�*:w'��l|3�_�[�g�:rX���`V"��l*���3�X���ۯ@Vk^ĳ��~b��4ھ@Gn��8�]/�6w}"��ԟ�ʩ���'<]Ӎ�l�8l9=��;Fc=�2w j�~u
��,H�B6�����K_ʩ���Xc'=_�@Dxp"Pi���܉��ˎ{��K��b�.�"���������n,�h��o�Eъ�� ��vMi+�1ʟ	���9��~��ȉ�5�I=;�;L���L&�~'���UcMѓ�H͜{w+��E�$���G�t��l����06�a��:�3`�����Ʈ�40������a4_���Z I�(�A6ZƑ��1�/��0�ИƔ��|��_w�n�d1�0I�E��hcS��ׅ|-�ʟYeE/�P�Y�M9��C��3�=���>������e�����x��-�dc��'T��Z��Րx\=��d9"���z�Y�;�R��Q�,GD��^Q9׀i;D�Qt�0�5�F�#����W��Y���W��R8���){\����S�z��K�z�
i�.F0���V�����n��x�I��As)��߫��7[26�?%�6g!���Y�A�D�OL�Fb�Yuy�2 F�
m-s1�����/�;�w��$sX�VOU�q�8�g���>L����ż4�II:L��c}kܻ��I��+S��藿��S�.D����md�lGf��>]0?�Rsl����L�T`a9!?���AװY��x�%j�A
s��:��g'&�'��2�s<�������讎��<@Xeھj��\:A�P^n\ނ�ݘ����D,Ml���{�������z���n�����B���ZB���9"lsh;#]�~��������^Ċ"/R^m_pQ<�C�wȏ�[c��5�[����������DDJ՟�3y���=r�h'PG^nx_��������/BǥA��M��b�t#�� �%}���6�E�����V��n`�'���:��K<����;�E���d�h��<��eX�*Y3��G/���mB��h��`5�U�h�D(p邕(���O}�C��T�jfɊ��ү+�I}���D�C�ޣ�`�j1l��U�	"�� 
�=O�QH��eѫ�`֥$9s�z5��VuE~��%�-n�խ������wȁ%����c�+_qAt��o� �m����"9�v`�<@
����!�hR4��H��qIz����0�g���6��%��?�wf�߄��Ӻ�=� ��� A��ů�I佚�&���˂,��.n�V��`�j,��h��m�����k+΋��%�.�ZJ�
v�x��q]�E&KBB��]S��4���
7�:n��ߣ����;��VSAY!�B/wTx���$[��:1k��Ł�DU���SX,��o�_|�j�/�T�6վ�p<���B��y��c�Y��~����uL|��;YХYy�Xn�T!2Lf����.���K����f�V|�s�A�[�B��L�x�4��t�dX������Z���4�%W����w� �f���<�O�o9Ԏ̟�5e�x@붼�>���=A�e\�h�pV��)`*�0�o�F��b�B���t��8C}v6n����=�?�{6���^��I`��ͪ��tM���",V��c����wY 0u��|+|��ց,�A�y�u����zkͫ=oU��5]//VWQ8�`)V��a[?���8�k&%F}�����!�l���㥎ڽ��7����I����P���Й�Θ�2=��"'g��Jkw,۫]��&CH)Q[�A���m���{��^�����C^���}ݵ��P`Vl��Wn�y�d,��L����������T�0�����_#��Ǟ�,�%`1�pU�T�YRآjO���� h���?(Y�������yc�\��YX4}����/>�^p��j��r����7^~nw���:��; ���V�,�0�@.#��|�ݐ�013X)]PY-ړ��xs�<���ݸ3z>^,hdz\-�o32��Ǖl�*���!<2�������F7�1m�F���]st���F�^�%-)��$�Lԥ��jQ9�I�ݙ{b���6gD�R��设$wӠ�b��X"��}5�g�W�fk-�V�#3�O1����L�ح�xz$Č\�]��b��BK �K��m�0�w�q� � ��O��*&�4\?Z7���y�����<�\8�g�n�w
U��V����r)�r��P[�=�14����
=�h9����G9�4Ϻ�`���r�Q�BQj�_��L�eٔhV9?��{ �0YU�n*��t:Q=�o��g���lDu��L���k�����<�ߒ�7�/���6p?�U��f4���`Ajʼ�X�]����?`d5��g9<�����7���y5�UI�{-��|R,Ψ�8����GJ]6����9�2�I���``�v�ی^ο�6a1{/���&��oB����LG�\͜�k��m'+Jp���v������Y/��c�k�k�'
[�F$��+:��p:4�@l�ޖ	�Լ�tt1`�ް�p?�q�/����f������,�t����Hv�-y��yJ��e7��թ�� �ɓ^�)����E$���]�����Q.�p�Rڷ�y��r�j����� Q8*'⻲s��7T���ZMM�dms��ԥ���$ș���q7(l��w�.�@���׻�`����D�[4xL�h��]L�У��{�F���u�w���H���u�����u��S�붿r
c"��o���$���a��鬱�u���`�˃1��M��f ���G�ۋ��B�"�C�|�+�qs��+k��ͼ܌x߂�w��
�ˤ�N:�(�zx�������iwW?.Z���]T�r�dx4\�����u���mz�]���ٙ����Q�BC�����?K��~��y^;��Z~:b��s��O.��d�ܾ�x��߯��{N�<m�6@2�AH� �=�y=���Oo���Dk,
N̐�:��}d�y�t�`�v�8��M�<�$�,[>����Ҥͭ�FV���$}�'~\�����ӊ�i������X�F����m�tؼ��IÇ����0�҇s_��9�4���q��]U�}J6qte�;�E�`sa��i7�mYp}S ޠH挺R�����I$��G�?>���1��D&��Ct����{W�^��ZF�Xۏ�hh:I�2��T.���tp �;ʸ$;n7��C�.��fֳJ)lBy�P8�\5s�"*'�Z.��_��A$��]��bm[L"Wv�t;�vu���L�������Qb�Ʌ�{�:���^��21��0� ��y#MD�}�e��ٚ� N����l�к?�����T�E���P�]L/8�:4z����l�l�Ʉ����((���͉��I���:5�>%�X�`3�>�.�%i����_O�K-�11���������{�3��Y#*�Ի��\j9�z�fWg�Q�7���U&�[�Y
*Hy-~��so�s��χ!]�2�z�>����I�s2�,��g�qÂl�o��F�>����8�=�aa���q5!��Q�����8���f�?�VA)X�闓}/{V���&�j��{mj��'a�U.N�����2���i�h��WSm؛A��i���J����7FN�@���
&}��w��w䊔#��:W1���=rNc�5�}`�G�f͞eR3�0_��ED�3_���������@D�T��퇫e�Tq���`�{�����A>�v=��k��ށ��Zf�VH8��B>6���ں���/���Q���ݡVy���=�[yS<�D�ZP� <{�-Y�/����d?j1�X��j�k���TL�s@|�m}qq�� ���j�Xg/��PHr�WƷַ�2;�鹖�=`���%r+�-ez�m"P54x*P� �QÏ������U�g�� ��+H�w�]u�B�:4�ٯ�ǟ6n<���5rRR��R7��J�c�XS�%%�'ٸ9�7���,/�)c�f���$$( �l��n]"�=o:úH��`L[>TY���C|���&���OԘ��RZu����"J�n�F�ÿ7�`��CA�<���]a�]\�9tԄ+>�|�`�pfc��	]��A:zǉ$2v8v/��k/l�p�'�D�?�lR|_8�_������P7�o��| ���	�����z���zdaK�DS ��W�u0�H�=wr28g̡�8Xj��+	�nT-4D���8v���E�,"8*X�	�9��}��t~\4d����2��Phrw�V�}#�g��ſ�.�us��f��o>򀿡���\\�&�R��b�����8��%n��kA�F�ZO_���7�FJ�v�h��[O]X��\��3(��O�o���eP��8J�����'�~�*.�{����� �$Q$��[�\?�e�zS�VK�w
��YV��؎��rYc8����Ԃ���?gʢg�|e��4���ER�m1�Ѭ���W{����8 a�.d1L�1�
��I ��3�MF�I8a��6%!<~ӄ*�&��l���ģ�n��U��M��j>��q��d�!��~���O�6�����1f"�oɁ=��ɴ�`Nda{���V��8ũUE~���s�X6ݹ=�4�m�����I�c��&:�
KwuՒKj�=`����j]��n�N�' 3YubyǼߘUm��$��`
Z��ɏ���K�G��,��U�`$�C�6Rk�eH��Q��<7��E�oz�qN���5l���3�6�����ډ�,-)��A��������'e�D���|M � ��a����VSs�A����>�N֖�/���'R6�FO�~��Ǽgy`��U���>��@�g�oz1� �q��a<9�a�v'|����GOXPܝ�Q����@��1�IΜ��c����
���cNڟ��;+	褄�MJn�3Y�2����r~�������+�R��>��`��{�	!��˸~�Z;ڭ]�	����<RZJ~�� .Y�!�=B-+h��x��֎W�J�b�168������n@�4ܨ�����N�3��7g��Dө���O�&��/X������.�
�E���ї�o���?�ү�0| ��l��ݜg@�{� �4/_���Z�0�J*ϳ�/���>�1��r:��[Pk~E���Nɸ��Ԑ�G4J6MU5��WC�\�ω���U~	��2�֟��J^%����ШT�?ljaѠ�w ��N\�E���6۴��OJvl�Cm���iҢ��W��
ɛZ��IRh۶��֟nTn��5�� �1�	b�|�kq����{��w����L�������|�.���_��4������Q�;�
�k>�[n��k�� d�-��>~�^�z�2��gƇ���UH�RR+_�b�ڇ0j�6@Qv�q�-�c�����#���8��[UĆ�
`귂!s�#S`#���[�Rn��_S��+�H��v�#b!w����o׾#�gt�������]����-7s������@��T}�,��bzI�G����ו[z�� s�U�ˇ��P2�5�Vs�hW����e�>8��c*�bci7�sgG�]m2C.��bi�U����ԔP��ɺ��Ŝ�]��+���K��5����9�����I���.�r�/f�1iǣ�i0O�i�+�ce���.z~�c��U��>��wZ!�ܑL�|�w����x8yb`u�r��a��}`D��p�%L�2Њ�ˋ�sj�����(��iñy�б�9��~�u�/� #��%WE2i��j�w�/}��"�*_�p��J�n��
�1�>k!@�v�(���>�a��&�;�wQa;����O�'u��
D��M�i|L�ꤗk��CL���t�& �;�$��� ㈖6W�i/�i��({G�]Z0�����_��v5v7Se{��bu#���r�[�%o��t�~��M�<��9���w�cb��g�W}�ϤYw\��i3�&���=0:����6���}'���bC���l�g��V�\�?�qC�r����S������ݘ=L�]�y�-y}n���_Y:���RQ���
F2����8�8~:g�i��r��A����ǧ,-'�f�Bh��I��=���k��[`�~�|H6��G7cFj� ����c�%dq��#Xc��.�=������_ ���� �zm<�9�n����,�N6����S�Nu���KKzv�J2���Ĝ�{��Ts4:3�),L������O���/�����aj�o2�9"���^������>����H��#�R+��]�i5a�k�b�����Q�Q�݆@mw-h���w��r��ӟ~���U3�0�e��<~_tO�{ C�~�_)�� 3o �R�G5�јN$�?/p /E�Y3-kC~��8���1d�l�xܠ:��_�}̧s ��c5�hIH���;�P8�j���y��Q������9��J3�����P��b����pS��%��Bv�'yo����  u�G��=uP%X�����#��Ƽ<N3JZ]��V#�@Ka7�����'��z\C���0��� M�޷�m��)$��DaϺ# V�';	  |������DJ�JI@��/&��o�j��j�T,��K���xƄ��?���|h���s��ˮ��K����7�T�Q1��P�VqP��+A	���n������V�@�U������If>��J���a���a��x�u~�w}�@�u���ԣ{xg�����t�_\�U�������%r���sTGc]M�7A6�u���c��.ԞcQ$uu���:Cmc�ʼxh���vM�su���p��`E*}3�Ak[hV�_�d�����&u�V����]�ov�?@�3d��W�n� �
(�5�̖�u�F�L�>�u�)�}���@۾�v?(P{?@Lv�)�i���Nw�0�;���$Z��U�ǜG��cO�`�����YK˨�{`�J��������:d���?���xG;�dP�����]�\�������oz-�h�#�{�)�B:ߥ�V�KO^�@g,�t���?�����/A�A�Vjb�'3�����t	��R�1�����c(�9?�.?���Zކ�'�{U�S������^�
�5��l4��U� T�ĺ5l��Q���[�]���2D�nyW<A3��J^��_17rf�O_���@����,�Ժ���D���XۖŦ8v*�hA��(���S��ʾrrէ���j�Ő�=�wqi��G�5����f(n}��ܕ
�t�[�P<xk�e����TY�b��eT��'�X
?_#�}ua�vWG���;0InYhǡ���Q�O#��{%���� �K-�@3���x%�m+�����Ղ�YbY6c�h���Rlً�JΥ�Q#a-W�1Xb����6�@�S:/7@�z��d��Q.;��I/�<������iW�W���e�! 1�j�H ���ᗡ{�'�nU >�ҐHLf-F��2��C
����]��3�Qs�C�c�n ���s�h�nw��*� i��IIYa9Ǜ�����8�}����Qwմ�Y[����N�T�ǔl��^4�os*8j{I�i6y�f�J�2�>c����%�Y!��������~z� ���5W�Z��{�jg�B�M�c\�N��!��qd�@��*�ul�����% �\��9�d�u;LS���4�J�o��L�6X��I��֒�t	K�ޚ����v��pnlO�:���$�}<��X��ٳ����^��#�Vb��W[�v���`fά��ث�8��4�B	��e-�u_�&�a��Nc�V�"��8��w��0�&�����I�;}I��a�J��1}=����]*��p�n����o��i���7)CŠ�U�bM`�� ����#���������q5ѡ:_F��,��z��O� 8{v�WO�qs���W�̆�����k3�>�GG��_��i���j !X<���9��A������d�δHY:J%,nU��cYk#(8殳kI�v. Ps�G,�N40�� �$���|�,B��������P�<-��lC����������?�J��;����}��u�l��%-������w%3�Y~cӆVXMA��e�Nw�zL�n]���{��O�6[�M:�Id*�v����)��Hvq���cz��e�֏�� D�ų�ߡ�+fS��(�
��%]&@]�����,�m�0�;r����+Y��{��ƃ��ONȿn�jo,�d���?��󂩕Udz�"�"r��9LW�$U�A�+�����ٌ�:���ߡ�8q1��:���%�R���=qӐ�0e�k�a4�l���[��솮�Fk(oU(���~�w��;���x��?�Au�Y����%�ٴ��Xzz���#�a:��û|h�"=���e���d���W�°�Լx�0�}LG�$��P.(Z����D�'T{�o�ܣ���܀g*��RP�5�2֗L���;��)�Y���ӊ�8b�RF�}���J0��	��h��[啨�Ͻ�{��Eq��3����h`wd��_���@꬟a�����d_]�$����n�n��ƙ�?M���=�L��|�H�٠WZ����Le��B\�*�m9>�*]q�J:�nl�D1�%C.ۘO���D@�k��\����jA^(U��� z���h����W�eY͜���/�f&߽��޼.^U&Ņ� OQ���T]���Q��2-Yj�Ļ�RW�WVe�&��������V�)t"�U�V��W�|-�FzZ���lV����}�3P��]���<����ס
���ր���&^/�R؋;J4�q��>���1�-tU9��y-͟f��B�
�Tv��V�z�/�K 0b'�������F�ҟl��6f�SA�F�� ����(7���s9��̀'Y坯BY�;^f�'#j����	۩�������*_cƋ��5�[�9jM����6t���-���F��1��`ʞ]I��/@�ٚ*��xKdSu�2=}��s,���_j��2,�:���Z����L�N�Џ�P�^m�mڍ�x�1�/]�4l��̍�zh�=�,�Ad���&�w�ܒu�������Eh��t]���Ը�__��3)g툷�1bU܋��G���0��<$i�ao�� ;��$�ۧeX�~Śf_����?(n/�(t�1BȲ�fu�6}��Tc�=��- N��?վ簯koi��y��HQ�4��a�j�y�c�t�X~�ϕ3��B��Fc�%��%�R�y`(��s6��g�"�Ƣ��VN�%��!D�GMpgک��uv�UQ���߄4JYՉ�'���Q 1�����F�ۀID��??��y�ެ|'��� 7F���V0�Sl,}G�mrb��$�u��>i˂�^Y��6�{����0�8��O(��Yd(9�����N>S��m��!,)��Y���k]�E!������{iC�l��l�2U��+�,L���vv�����S��%�*}ߍ6�s��PL�w�x��IC@��8�tx����sڹ��<��ޖ�����,Z���Le��ܲ�V��S7
�<./9�_K@MSb;Y3�F�F�[d�@��9�Y�ᗁL��&ƨ��͗7C����S�����7<ng�\p͉����ۢ͒��s�`�\^��%&�=ޗT��&�ip(�ߜ��a��%�kw��cҎ�e\�8��l���s��e�Ia7��tJ^������wIEъ��I��Z��~���6neH�B0��嫹6�tޏrrf�[�A�-_M>�M� $b��O��Mr\{8)��3�@��{��ʐA���Ŋ�?t���xz}��6� �|-����m"��NqT�:w})����\��-�c�7���=^�ZS5K9�]�X{����e����$��g�i�u]�Q󳞁�I�>zҧ��vh������qQ$��𸸀Jr Q�]�$Q�� �"� 9���s�AQPI*9�䌒3��"Ir�4�0�a~U=��|�������Uu�9�[��7� ׼���嘪�Pg%�����\��m����n�-�{���/�������"N����S�����,�ŉ��J�D��Q��`�E��@9�Ԑi��A-�$r�O���te��j��dEհ;�&Eu�5ܕ�ӏ4=�G(��(�+�cx���b
��y޿/�5Y������-�ݻ{Ms͑,X���O�p��?Ű���&����T+����s'	��wq�t�Ě�6C��0��N�2i����)�O��p��1��$��JE7g�mѲ����GqVI���Be=(��������-�k3`ť��Ӌ�7'�����*��J��\�K�9*������W:�R��O#]TvJ9��n�+ˀ�D�B���g��K'�nE�<2&U���h�J����DM}jsŃ��m�R(� R���Toh�����^F�s�;A�b3�n_Z@��
�&R��NͩX�tpM%��S��DP�V�zp�k��B����C@�M]~�X\������p����ƙU��ߚ��\T�g+W�x�����#��Ovg?��_�r���?bǕhjy��SE�?�#Ҿ��ʞ����q�������fU<���y?ٹ��#����YO�럊ˬ��!�wh:cgy�V�;�c��:?�R��n�!�e��l�Ad<�0ǃ�<��Q��*�7�jno��
�T�Avd��������>���X��rr�ZN�0��xF��u2���L��{�3�U�5��kBEsobBf�3gC6�s$@�8��&�Y!/���'G���O��WGG `���[x$^����*�����E���E����)�M��Ծ�ۼ3��@g��l����Q��!�:zb�B! ��%��!���tw'Qe�!]j�Z�"��*|��'��:U91mC�zu�e=h���1�<Ms����˟QF��]oDX�R�Cޥ�e�����$2V~���x5j���<#7s�UÚMT��T+���)6���5X�:(H�ฎ��*7���!ۏTn�*�{��p���������D
!oр^�:s�/��a�P.L�j�uX����ޗ��w���_��C�w_�n^��Y��	����%�r��х��@�6l���(�T�,�R�h�y@�}���g�.B���'�ծF���%k������xo<��O-�ziP��:������z��ӝOa�"�^To�*RNqd}烮��nX<`}�O��3k���QJyp���ȇ�S�&z�X���d(����wǚ^�@CD���6t���$nӛ{89�w��acz�:zN�X��s�|� �v�1�,$9�dY��k���0�O���Q-<9��qw�X�R<E�$�h�W6ܮ��|e��ˑ��ٔ�瀼t��J�2GL�-��T�	���ʭ�$�+e�*u5;��R�7��vܕOfwd�������:$l���Kc%h�+�@G��]���1�����cp� K�	��K>>'3?U��YleS���Q7��a��ٵPk�Y��^4�/�B�{Ng����;�����q�MSٱ6b��1u��f��m��Dt���f��;!�x-i���ܽx�}���g�'�6'z�)�_/�4z�	~��2�i���`wP�r��BY;G�v=���3FO��7�D����&�g�R?��j�|_B��@AN�0��xP��Ձ����β�d�$�5�{#Z�n*Q�cԯO��8i���ʍ@n�p��[\��'>l5�ӥM��,
8��b�Sӛ"@cd�^�8���|�H��#�RLfn����5%�^�v�]ﾏ�2���N��[si��^��J�@|�wծ{5�BƨREm-�^A�R,v��_
�GNS�������8��_�v�&��-OM/z��w������o��A��Jޯ��P���G��/�X.dZ����ֶYD1��τ3;	nP.E�d͵���@������v#�=K��e�(���nފ�A�ɹ�z�y[^�H��gs���|�+���z�[ӣ;��d���7��]�I���a[�S�7�R��a��H��'�)�����N��[��tu���.�vegg"����!���O�Z*I�zގs��`p
ܡUv�J6",��κW=�6�c&��p�����Ҫ,첥���m��9�NVҸJ��� r��.Zx��!�����{8x�Wu��PQ��%/`�VV�%��"T��N�'�7ÌR[n�|������~
�{uS)�vU�y��Kp�8�b	[L�vp��A��X/����	9�m��i�Z����\�L��t�����ˡ�"z{O�ijp����.E���(T �,y'���rv@|���a'/�Gߏ8Qc�	{g��n������̎�*/v���Ce����$l(O�~��<�O����x�Su�
V��)�+���������� �JN�ɖ~�6�B��5�G���8�!yC�f��SQ�h(Z�T����-;�j9��7�l{3����*�Ϯ�>�q�ZB^�AQ��l���	L���ލ�ao��H�!oB�Y�t�JhoV����넕��q��ZbHk`H����09���~hz�d����$�>}��k�"�W2�> ��M�2�6L���qǤe��G�6=�y��}{Z1ٵ1��b����Ĳy>���쐓���wqq����f����c,!C��5�.��e-������<�+Y��dl�^z��892��KiE���6@g���Wfm*/X�H;�����
 �3�'�;�C6�������If����Ip�R����fa�ލ�����s�#�
�I��(�Xi�����_�eQ��"���ٍ�Y4�"�{�$�����3t5e���l�ӄ�dB�r��'|>�2܇��tZO����vUR*��I���͛� ���M�uq[$�yQ����k?x̋���bzGdA|�16Eԉ�M��3iQ����� ��_�硛]L����ʙu��B�ԟ[���]�����_�%ZI�U&|p]�b����<ؿ�3t��!�}��-�&��_�lǻ�:�.���RN�+���H��U��$Nu<���n	]M"xo������F��g-�������.�/l`�k9�ްz
��|3�9@�ft��r,"g�����w-�(�\d��|�hz����o������HU��T����[�u�i0��-;��p)�ߦ,������{K:��)^fh;7�>pTLE�a��>cR����>jԙ+�O��5XK�q`&�����9����?�^Y�8t���e���v��Cр������x�\�Ârl��G�H��C7��{�})A�y�Nթ�`S�ޭc���ǧ�V�;�3Ww��g��IH�P��/U���?��pNNn�m��+`:��芋��(�|�qʄ*�TS&$c��l�-6����2�>��vܪ��E|�`ٜ���i�2t�g��=|_CFT��7����F����l��c�/���|�O�����r*d���@�~��
dԍ�����h���̬���t�����3@�z�g�1�7�d�&�"o	Q�����v�=T����]U&�CMG)n��͆g���,����k@л,���M҇§ʍ ��+��o�L"�3������5 ���mn���!k�Ec�v�fV�4���/3�J7S7�~X�]h���?�Zj���Ju�n�:�R�6)��/'�mʲe��8��R�5�����O��U�%Z����~�RMW[�k�����n
ɝ���P�i��k��'Y��B������h�2���vhZ!�9�`lcq��9v�Z�V���~{����F͛k���8|�0��]��H*f��W���4t�+��	�;7I�{ER��ꛗ�R5���&-�����e�~ys�ڭ��P�U��M�e�I��V���}I�N�ѱ�KT�7j�Tc�%�w&:�ʨ!��8�#%:�����E<���_i�\8|-�@q7/v �$K�sI*3�?��2k�iP�T�m�BXO�njj|�-�?�z��.�7��Wa�i�so�u�n��@���`o��!9� Kl�=��ul/5吾���}��`v�^OK�ow$�ߕ�%�1qϛ���8��/_�7��7�^�L��x��΅{��zɖ�O�7�P\]s��u�V���;O4�z�%��fs��5[U#`��IĹ�Rzn�]R���a:����؝���9,M�j��i�Լ�P���t�e�˕���Eh���_κ_r���iZ?�4W�S���-3=�$dq�<3@���ΎӅ
�d�OG>��Z�&�:�z�+p�o��5�X���/Z%-z=q?��nq����DZ��B7�����G֙�6e+�@���j�z196��"P�B�����wm�a/�g3̮����g9�y��#.?3lrr^>��f���o �fWlDp��+����h�����L�%�n��:��%aNE	������j�(�D#������y$�1`"���7 ���>~�����)6�bnBo��/������bo!~��F�@7��z�wb�]�ٷ�ub����E��m�^lR'�,)�lr�� P�N7*b}�]�������[�	�E8 |�RL�,L���Q�,�bl��d�I����2å9�˲u4��� �-��C薕�p� ���r�1�}ʆ����ɢ���s�B��V�	���A$�$�q1����z1/ďQ��g ��h&H�ϐ�{����
��L�^D3����<��wǘw��e&��@v7aB�x��m��s���D���ٻ�O^�|[d�!�Z2|7BD;����V��|3\��#�F%'�u�8-k`]�e��ߕ�.>8��aN��1���xW�}7����*6�
U�P)�s*�1��58�+����ŨSŖ���QF"G٭<r	V��2#s��)ݰ�����[L��s�3��?����������m��!Q�h�$�r����<�������sT7���5��Ow�I|Ş�s�L%�w⣖���T��cf�x�3��+�<~_UZ)�_�/�zt�b���|�X���tѯ�i�h9���n����0������>��v���,�\�g���h�qT�mwo����=3��^�3��c��/Z�mS�mk��Ź��z����9=\c��+�q��
$4���Z� �ɭ�0�>�4� ,��)�Z-��@yv��|�n荎���4`�"�,�ħ��tɸ���Ġ�����M."��m����m��}��f2��o��>����P�g�鬪�.-z��t��~ΞO�Y�)��sH�x������d��T�<�x@�^Ui|�V��	ź�ȗFQ���3�t�@��ނYk���}[z(���k���M�zw�3�B��r�j�ܧ;�lw���sY�!N}ƭxʮV�R��:����e�Ta̻V��e��.i|�p#����s �f�dd��*&w�!Mg���l����}��T<��:d�%x?d�K�.��8/7��|��g}��g�\�6��Xq]K�5i��7T0�Ҟ+t�`Q�m�9����g3�� Y���n���A���{J>).���i�7ދ���C�;V�>X� v������Z�D[) q���w<�wy��52�]wf~����;��qVg�t��Z_�$����k�V[��1u�@�H�y���c+�����Ob��%B�wg�jΈ|UtY��t��D({=�	V���P�?k������u������1�X�[	���W3��
�O�<����4QRƵ�e�R@}�>�&��c7����X/
�H�*��C)F��Ύ�Lc��l�y>��"�n����t�a%\����x���ݮ�ݻ��5�Q�7�ݽ��<�}apf���>^��>����'/��s�|%��2O�߄[Xrd�a�7���K �I�;�`��y���x	���r�<M�p��2պЄGiP<�PP��T�Xj������Z�9�Vw��=J�y]��y-V�*����ur_�8)2���b7�D����\O��̹�w���PV�3�?#�bq�
X:��-����Q�ﻗŭ�ϚBݤ׃/.w�ݓ���e�1j�)X����vu�I�5%~�l�@���I��?��5t�j|@بa�8�@A�0��Jش�Vl ~�5���.���C�F��>�`-��Y�eߟn�cpf��>X&a��i��Ic�^�Y�]��T@=���	'�<����P;_x�L��lh8͋o����k�����Yj��e.�x���q��բ���& V��9�<hI�����M6�������i0�o���E�[8����=O��cz��C����v��j�"]O�<5
�\��(��B���dOJ�
4�0r�~�0i�����xi�C%^�U9>��/�^�Y��kٺ��H�%�A�)zuw[�C=�7`�=��;�eP=ja/�G�Ul��T"�iR��c
��TV���r�g%��s!��p�%�t0��d$��°�����-�d�*�������=��uu�H�&��P?w�t��6�kT�?@��R�vDH�{������8���9��冷�:m\(�@�?4�--�љ:Gg��ۍY�Q ���|��e�%ȮY�$%7K5�Q��Ke����ʙ���v< ;�ɸ�'�{s�!�P`����Ϋ��C�^�Ul�ԔO����2���*R�:���"����o@J�����Gg�n�U�Z4�%�v�жLͽ�O�SN�~ҡ��b��\r��ʈt��n�����d�UX���&�NX���w��T��b2T�X�Q?R�"�J9{AL^}�@�nfo���'/�σ�MM���/D�]G�qV�{��������\9�3��g ���U��gs(��Q��	X؈�k^tM����K�a:[`}\�c"p�^.�b��(%&ġЪu
��nO�7a��u�Z:�[mR�$�F���軄蝚��f�� ���:g;��	���P�]�J��z��橽-��_nSX��0��%P�,
'��پ�K��#�ًE��Bx"�"`X�(���?
����wy͞��%�[��fQ��I����n�nX�G�#�&/�?�n�=����#t[˔���U�M�AY�c@�+��U(B��P�d�t�g7��LC�����TvY�!��B�SҘ�F@��}���5�o��\�͘y�P�D�� Ƿ�`��+�[7|~$�NXظ;�߲� �*�G�>z ����("��.�k؉p��-����*���t����ށC�v<ē6TC��s'�IND xѠ����h�q �WI9�y�ݦ�E_P��l�U�i�Z���&;�(�"X@F3F�I�s�2����ݕC}{�.yu��"�ɍz}}�<q���s�֫L7��n�P�����s�W�5�R������^�ON6���B��1'�U2ӻ���-,�����^�7d�$�R9�w��{|�9!Sro��/z�H�Vi��E�*�ȣTf�d�<���� <@`�I��?ΰs�>�f'�
������v"E��D,�)|mU�����T��S��]rG,����7�e�N�d�,���EK�;�����-ܑ)��q�/�_ƛ�a(fŷ���4��g��҇?&-�b��$!}�Y�����!�	E�@j! ��٣LۊB���FJ��$�:(5D��lm�ƍ�X���bĘ�N���b@8��>�d{��!�^-W��!9��i1���ы�C�)�^B��}�:}P�
��X�+�J��.ƹ_d�D�/��{`����֙����	�.ŴIh�ZD>j*�����7-��$:đ_l6،X� �S�R�N)��	��{m���}�Hbaьߣ�-��ߪYF/��Lah�(�>iH�R椂��x�����5I"��.;P����r�e~�%`�i�~��4	����R�k*+�&��~g�_w�@��%���p��c ���lZ��K���{�Dgl��q႕C� �T`��^�����@E��,7�\��o]g>�K�?fF�8��2g�]h�`��{,��P��:8h��ijzZ�	���=.�v�5�	�E(T�C���j�MqZ��j��̞7�4�X��P����ooX٬�;�IA���M7��g���O��'��4(]�14�h� 9,�ssT��;I6j͢M���IN��kL!��2HTJ�1g�l��ʋ��kb2�K��ސ�[w�])R�d-�J���-��uޮ�"w�;�c�:��[��:��%��ݭ���D������I�<�F�)NՆ��EJ���(�����X���|�]J����i��Dr	։;��ðc�YS�P%|��әX�Oi��������������F�1U�|fծA�H&}{�eF��9��� �i��(��s���4�ޯH����[_��/B��9S�Oʲ[��8�E+�$�IH�N�u��lnW����*#���pΖ��6�K�����#�ࣦĀ��v*ƽJ�e�<Hz�����"qmw^�� .9���ΦU�m ���a�n?�| ���o4ܾ߲��d2�Ñ��qc�eb�~ā�I���XQFl�qB� 
5������8�^n�~�Z��"�*2�%��a�*��ׯ�����zG9��rj�dA�I����j�ì���ү��?㴺�H�d��rl��!�@^�}�ZL��a9�B�n�������, Q[�S?�>�P�Pc �f�>���N#z�$݄H��L�|�	��?���,m�[;.u�b[���ٸTߠ��I�,(��]3AҾq��NW-PTh��e��ϱ&��ND͔Џo��ޖ"�B�b�WF\�1X����u>���/ƹ�k��R��M�,�c���[�p܌e�]���¬���y�U����sX����|��T���G��*U)&N�*���,fFG����X�|_h��� O���l���qGD�x�U��X�
�6�u���t-O.�c<L��)�@k�������S�k�j�Lv�CC��j�uN�BU<�$�/�����`]��DܷVLC��9[0�h�;2���g��l��5�@�NO/.^N�D=~��t6�dO��0Cߗ��R0�����/��! w��i@��d�
z��b�j�z.?�A;��%�l���ޯ��aV�}Чښ }�Grُߍ}}�,8�=m��=��K����no]�\[�>"�lw?]d�о�ߨ�:E�\8�$s�p����<ii:K��^ �������3'����o�p���D�}�)?�|9��'^�d�1X�[x��Oo��R{��@#����7)��8�D�t����i�d�	����2v[�ݩ��=����R7��Q޿�Wxn����򽟢�QӍ�P���V�S2�P��H�G��J=	]��i5{��!l
�x�$pu�7�䊘iE��n��M_-!3xGL�{��6{x�~�����s����MmeP�ɤ�n�6����k!�X��JfEd&����k�2� ��
����٥��C).۔�����?��خ�#T����I�E�&w7�H�
�i��:�����o,X��`�\H�9�'S��$��
p-04���j$
��ݚ�f{P�E���W�{:�w���F ��#Ce�M��0�^�8�~�p�F��)_E�S�H��t���ws���R쎭�������X:���vPyoM~���XR�Mҡ�޺���uFF�V��D�ѯk��Ѳy�~J����.]��.�S�s8�hɃ��ǲu]g�"*kw&�s���!�E��| Lt�Z��<� ��Ώ�FEm����c���_�M���|������z�#(Æ��'��jݐ޲�]K�e��i��<�C��h�h���X �+D�V`i?���:~ �O��*���7��V�v8-�煮2$���ݟ��L�� h�x�$J,.��4�"7�mȻ��D�?5�Q���HSr��T B�ݣ6�X��	:΂�5}���`!s��v gʤm�m�����L!�\������7J��o�X\�b��2�L�bi�%R�Z��f�^�/�D��jTL��>��S5d;���|��G��ES޸�D���J�۷�)�P���%�bI�p>�`մک�
#��I�8	�	�ЄQ��OJ�Y�,�/�4�
��f%�k��y�Z/��A�O�'~}��8��ڸ��
B�G��}T���~Ҹ(��FJ���5xx;g,@� ?����T�=�q��n�1z&"�#Ч1P��W>M�/�P�Ӱ�)�3-H�G�uf��)<�c{
Ghf:��ȿi��ٶ���K�:O��Y��'�)Dq�0N�=�E�?	�%��D�؟�����h5�xBj��	�*[T������XS���{�(���j ���}���sp�WM��� ��<�����t+��)`�I����1��|̧##�ܬ�����|�$2oI�L���L=Bg*@̮�q�O�Ty��*_(9=g/d_?�E;�/��LZ�����z��LH�]p�^v#>�2o�`�x�Fo��hD�ڴ�?F�m�v�%���"���7�s�
DJ��W�f��~�FR���$o�J$�7B�D�Q����*@�%�g	f8��w�`�1h���TNf�.��[� ~��ӡ�� �J��<��0R0�bS�z
7���n��e&$t�T�Oӄ��P���3-*pb��En�ju�t$$0f�M�I�mS��3�3���-D����2�t�p ��t���9�v�@U��9̯ˮ�%Bd� �M�!a�4��P'�ר���s���9> }	*���E3"LO��(g8]܅���������2l����!�5^�Ϝ��R{y��s����Nɖ^�M�t@q���Ĺ�d#�T��ƻ�c���0�obBჯ�~{�����.;Ӡ�;2O,l�ʐ����������"�xc]')�U�cu�,��bت�v���gia��>&ٳ@�����a�AB��}.�'��p}.fg>�3L���O�u���/ �&��;ޞ��V���q��U�f��-my���$t���b�3��t7�j��#����M����&!����1Н�TV��1����K�`7�=��T>L���9t��'e
���B��A���2���Pv>����I�,`�� #2�D����#�z���&�^�-]��|����O����gu��ch%�.��1�\]�$�\�e�ZN���υ�q���ۻ�d�*�n<m�1Q"Q�#��u5_K����:3!��Uy}eO	�ӯ5 xՁ�M����=]1�9j�@n%$�M]��ɽG����7�&1a�Qg&�x�%�.F�NRu4�yqI�\3�c�-� ��t��6�`ǫ�
0�ÿ���n6a�b�@}$W�W�f�AY�$��N 	��CJ"��/5���
���!MSѻ�W!�� @�F��:��|�[���|2զ�6f���]r���i�D�'w��fe�K�����^��-�!�βȁ B�\��*r�ut�fZ� �b���ں4*���(j<��N��P�&g r�JT[���g�����B>����tk�L����>Zo����0Cݓ�. ��-��`a(4�����T�C�Sg#_�6�e2i%��t�Q
��haS�Z�G1�5_Gr9�k��+==�O��]'l6�@�o�ıN��i�ݍ��1�m���8b�P ǩ�����
ÿ�O���`�����`H�Q��&���~�*�;���O�8H:ȁ�7_�~�+���8̆:�!'���Y�q��t�dT^���+<yk��Q`���=�v~��Ab�U��}���A�6���RlbH�{��=���ٱB�J&����ן'�v�9A÷��,�� ��~�z'p7gw���h��\)�7k��+��'���%��J�	�|�L���6�9�� O���~ޝ(JG�El	Xr���QYP�a�R.��#ϸq��D�h�mk���7��R�]�Ӓ[*�7ϑD��R[@���1�F`����9Ӎb1q�"�F$8<��
]
���EU!o����8�w���UN��i���8����Ɩ駞�M����+����:yP�4�����UX��1gŋ��_ix\haU���X9� ��z@3�޼H?���c �M��GAz,FM�KDBP�9T�w��8!J�jf(e��
:��u�XRrS�I'@��۔�6$鐇5�a�k`7����o�tmJ*Qd�u�b�EdKB`K=���` ��wY�����Tp[��;(b*����{'k��	��L�B����"|^G��.��
�C���Z����&��;PVVI�%��?ݶ���yaf�"DU�Q/�84aX�Ab��E�����yE�@��Fd��A�	����"�bl;K���b|�'�6�	h\��E�@��Xd~�\b�Yk�����z�,6��~Ŏ�柃 ��m"
�
�;���y���`� ��ʆi����K�D�"f�k��}��Od���a�9Q9��P�X������{$�O.�,����k�j
M#���(@�_�R���>����a܃V�������O2��	�͡����] �� ��Z�rXʿm�.a��DiN�e�v��anԑ��M\&��|`Q{_�*p�`���'Y�+��-�H�f�Ɠ�uC�II�� (G=�<�0%�/�j��f��e�������P^cc��_�V�{�.:�G�n~��Zq�8��?����re��%`�5D��`A�s�f��O�cAfE� e���f�9P�᣽3�5߀Vq�ƾ��4�EϺ��������D�]��;M`F�n@>0ǂf�4|�o]��*�2�L$��ɽ�rr4�>&{Q��_�qp6�y�`��D�F�~�NGJ:�E%$m�.��F���2_>�+	͟L�o��qU�J���D�h�2;z"��� �7�L��z|�G+�6�������x��D)%��b�I���Y
��o�'�������ƒ{��或/3� r	1U�h 2���=�7��=�Gu"��(so��J&���\|8a��������=�J�
2�w�)�j�`��\�Q[R@�`S|B4�����
�k��]��%��2��K4E� ��}�6K�F�J:M����>���k�6b<H�̩d��3Rg�����I���$]4�?'m���Ue	�Z}-����Q2?��cD��R������a����:I�-�֕����^��P�~`�V6"-N��ȸ�e�&�T6�t�
��%��vւ�i�`���xݾK��/K/���X���1������w"
���G��0�|�p��p��7g)�T{�\i�G�Ư�bc����8��Ѷ>bS�qc��!����_�=���s.٣©�*:�zK�"�ܽ�׋�o��elOq�������ҡ�򪝎\F�X"[�Tg�?B���pa6�2�b���Ŭrmn�O�
��Z��qHオ���',`�{?�0��]H[�:}dҿ�[��������9wu����wJy�8��=H�5�z��-h���=�3h�A���;ҽ�]DN��?	P���6l�[��a�;�xKɒGG�
��>9>th�yot!�T�`P`^��#{2����.P��n}8G���̌+�����MzW��9�4?�;K{�-�g$��+�y[!�Has���E||�_D�B�<o�I��C3.{���4b'��,�8��8Y]�|ʑ���~~���j��Ü�x�����0��Wh�xө��`IdXslL��v��t��Xn�j���Aȷ��=Db	o�ֽy�G��՘+��	a��DD^��1��W����~�3E��4���--[��X��bQ��u�����&��U�H{a23�
�P9��4S��i^�v�R�/dO�|#\�$�V{U����i�i4H��Q��hGS��@���<T}7%2=�eq� F�N�W�6�p�0u���+���og���pu�B,g���O������ XK��L�d�]�i�8�b�F��+Mu�W�6`��h�֯�Y�!_��\>�͝���I��o��Al�_PI��xK���3퇂;
�� ���z�Ņ����G:2�H��d.z�D�4 ��W�
2�̭�S���z�e��Ce�����1h��q��ۍ��u9�N����N�������+��o��`#�m��3P֍eNI�`*��䊾09C�U��ŷ ��u�2[�f�l�3���[x�ԃp=���{�.�e׵-�|���Y�!��e����]�'���=:�`:���5����k��V:�5{���*F���t-`��eaY�*n"��"jkw*�Cֿ��^�d�<A�Hw�&)*}�_.^�j��PD���c� �hj��?�F�܄ݱ��S4wʤ�k�m���<��r,���>J�ƀ�����:5��؂��:��}%��Q��r�ޱ-�cNB����6��_����b�O����&,%�fl?�v|e=c'(j�^k5%���DϬ�ܣC�r�M���!#L���z�3��a��a��!`�m�L�R��v�l[hZ�ÌB	y���vwC��(�����=�.i{���v\!W����u9��jPX�cw�OY�w'��}��V���#� ��;۵3��J���ɤ�T�M6�mA�F�ֵߗ�v@�I-�f��b�2����z���M!Z������y��Z�1X�`K(�Z�0�@�w��-V��d)�<H�ӧ�(ں�v����'{Oמ�Z�n��1��V�a3�#�l�;{��kO>oѳ-���;}enh`���Ə�1��k���K�t@Q ��sx�~���C(�`k��
ZS�k� �$d8��S\4�J
{���=q���Au�L�X�]�$��þ_���44Jy�a^��b�IQ�-\��&����RnP�eNh0�~��RH6I�x+U��b�\*�@��K�9��!I5�o����R(v�J:)��\�v_g��Kh,$��R��+O"[����#�`j[E,
}3;IE� 7�*�6S�i��]���
��W;�N��R[U�lQU�_���8T��pngq�:]KD���"�?z�6.kW��T��&q�אۻ��.=�4n�C~�)
��DB?VU�n�m$G"��u�2=�LQV�gh�N �g�B<�����ˇ��9�z̭;!*���SvIp�V��Is}��g�.�nJ����U�F�`�<㞢sU�����)�S�(u'�c�H��A�K�h�B8*	j�z�	z�
'���u��
�ỵ�V�:�DI������p�'���s8�b@��	v�u�ťKҚ����V������=C�-e��N�-���}<F���-�>4tp��-`�[n8�c��_M�	v2;y�D�,-b���)2Uz�rn_K@8
t_R\�_��8���+�`��`&1]����g,D���o�<��%Q�9�%7�%Go��$3zk�c��奊Y�R�� ���I]N�H�M@��זn�_K��{Ҭ�/����[0��;�G�-m�~%�P���J;Sݟo�wP)u8ϥ�z��l��0ɜT�`}?�FUG�8�=�\Г��C�~3���>纁�a#�Dyu�e7���d���j��\=Tf�&��K�SZ�Ɏ`���a�"��P��'45A%Yۘp��Bo��N�f
��ն�^%[����wk@���Y����q��ѥ'e;��^��6]jq�g{ 8���‐S�&��%�5	��fʌ�X�d�������UK��CI4�îvẀ�	%lKݯP��D-P��Wf����GZ�˖%�=g��%�-��Xr{�^hK�VI͇����G-I+�_��8�Pj�0t�~ �m^�D䱯.�?�XN�U	��'��i4g��Q���c��j���ޔH=��]��^5D\�A�K@s
��-�n@^��
�2�[�:9snu!8�T���(�����H?H�v37P�a�{�3���z�*StT� "훽8'H���:�mqE�^j*{l��&�'���a4�A���7^^I�����`멜S>����f{��{�٘v�ZZ�Ǎq��L^ۮ��g?��I9�i9 ������o�om��`G��\�������b3�)q��u«NBP�:�d�6 Zo�*%���wڤ�&��&���ý�8�j�+wl����N$<�%����-/J��"��}��'�g��Y��~����!�$3�k����u�5&�t`�&��V �z���\����~
X�B��Pv@p���N��lS����.�k�\X2��U̫h��5�~�|?��o��7�b�^)c?oX�W��}�G<�U, ��l� �;�����$���Í�0��*7���;�L�9��N���t8��w��^M�����Y���]�f���z�AS��֑���W�b}��� (��@�:��La<c ���vo�a���i��L|�Ui�1c�`r9�1�5el[�I�s�a�U"���#w
�qP��
��6�2��du?h�S�A�
w���� ,����MtH`�; t�K���D<���3���׊��N0�-O��$��\fwH��P�B�'�Ã�f
���P+Y����s������-Q�K���@y���(�!H��L��uA�|�NuŦ���p_�rX	��U��n	�� ��WP&����m�@�a�������@�;W_,�zt�7��7������a���O����;�% r�O���Ђ��\���,�G��4^c/
�R�-S�� \J��vY�i�$P�Z�w�N��S|�BTD>mP���pT���\</���M
��qD%ᮬg�C�s�Ⲫ5=�n��u��E��M�M��g�M���v��b��x�2s�M�}�
��vGi�KRa}����;���M�G�Ѿ�<��Wjȸu�� t?h$�;πK��)�g�_!���=^Y���ֳ;B.�Ly����7�����f� ⍭)�����D�w݁���k�� �ۺ/Ht|^oC�t���򕌻{��{�VZ�~�e�)06w��z������fD�)�ϑ&�B*���x�#����������uW�4�mP����h�ڈʔՍ�������O��1?�@��m�����Oqۣg7:T)��������K
��ʮp�ܚ1O���M,���˹��Dn.���!]W�Ө�G%���:,��Jl]d"��Q����<���j��B�<��`x�PZV��f�� �IW�����ӂƵ������zt뿤�%}�uS{���Z?�݈NRQ�H�����b��&�W��Tb���|�dܭ�;�;�qU,�VPK�^������S'@�֎J�%�l����/�m bbQw�넧�ϭ�~ᇽ�-���X�_T�Ӵ�i$��RǛXLд����,Qx2z��-^��?����_���Uۍ�h$��.�I:js-?:>Ls�J�y�h��+x��6q��b�?�K��$�
ťTk��\R��:P��č�pX~��V����f�D��F=<H2�ۅH�L5=���n9f�eS��B76s��i�-��X��[B�����bs���u�x�c��nm�,����V�]����영Nb��1�ZŃ}9��ڟG 󵚥���0ԩぴy&����?k&1��?U�}����Z_��v�������L��'�嬔dHf3>nv�^%�Md�2�2}��4��p9�x/��q�eg1Ym�YX�=2����qb܏%��*�KCCu�&�9쏉�� �ۤrG�H�+���-�(}w㒪��Ĳ���Q	v`ij[^�g]�� d�y�o&�����ub�W)�%J���2s����)z��s�*�S0��W�<3�����\`Kw��q�J\F����]�o�ג���Yų��뻇��w]l�~7ch���$\cB��W@A	��K��f�3��r���yKMR��=�Zu�E��v�C��{��幞���>;�X-*��Hz*��r'�o���287��g顿�����p[��IM�+�!�;#i�%��,E��I�����j���s�6�w�;�{,��}�������?�e-�y�n�dp���#�Թ��jb�OW����w`-Q�j[	�S�e)��Ph��s�A�s�W���z������u����\a�ҙ��K+�J$y��M�~E���'�`����3��Y5�լ+�w��;1�� $�ق�p�]���ݽ��fC\#���Ϲ
(���+Tևڥ�w���'/a���iR����]���V<P���{?�7+��aVs�׼�$}����Yw�m=a<�L|���>���*(�g��<d���^k܄��{-llE�U>�GLR�� z%9;P'z�G�YF�S�n[#�d����]��׍V��`Q&�[}[����s����9i�Ѷ=f핽����4�q��������33�xC��Ps���o�ՎZi�حng�q�d+�&ƀ����LU��]����d�T��!�)��fef~R3X���-TGo��8�=ʇT�G��tn��O-x�B�r|�m'���DHٔifpG�rf�Í�π5�qv{I�!J�9T��KE�\��+�k+Ʃ��O%+b�
���q[�r�xB�\z�_π��1�T>+U�D�� ���J���i���Nm�jo��m?Iqg�, O\���ki��!�~j#�>0A}��u.�|��ĝsS��T���	�;Ol���I�/0燛��E������x��7�so��[��VTJJ��P2��m�PIȘB�1dO?E7�.�2V�̉�1���J(2�$�1�޵�^�{?���������g}���}�����*_�� 3���v'�˘�Ï@��}}1�����[o	w�ybG>
�+��z���2FTCދ0c�����6>{� s;|�{d���*+]�ٝH�]��<i0E���~��F��Č����fOl;�����%�ڿ13,�㬿�(.MƖ ���>KH���0ad�J%����B�녧�~ �o}k�7�_;-r��O�nJ��b�v��`����|�P`:a,� �x��Ir4��,Y����%Z�N}}��B��r�O7 X�Z����IL,#X4���6|��U��f��	�7��iH2$�lqX��K�"��%�STJ���T�+�뛋ϸ���V;b-���%�j�~t(,�B�������v	Pw)�BUװ��i�S�!�Yl�;����e���R4�G�s����R&���A��)�"S\�	�;��T����mT@Hqi�y�ga��:��&��,�z�
�zJ^���{tF�
<�?��"��/gO����w��xU�Y��#�bi����^�84�+����~Ք}(�O���@���ҹ�͏bJ�re�UJ/�q��8��w�H5 c%�8��	�u44��Xu��!#\QRH�8٣�̕Zc��S%��|�ٗg	��p�p=��1��롊J2�}�Gkp�N���O3�l�T�ʴ<'<Ɩ��6$��'x�pUZ�<���Aȹ�|�f�����E��s2k�H�R#@R��A��S���ւ��[��\��Kq$���)�����xH�uvV֠U)b����k�7r��[ ��S�>1렔}�ίn�8���= ��U0$�w����"���*7� t��v���O* .��7��N�8g,��7R��̯?�A���c	t �"u^\U�ʲ׽��w&�rIي��^O�[��m��.�j0�V�m���圣���,�7�4~8��~RS��'A�tv)�J�; �Ȉ}�>Tx���{�z���p�n�b2������V)��V)8L�m[eoo�G��KJD�?�v��5?��˫�I?��R|�#�����Τ�?i����+#�{)�t��/L%<8C��Ɲ�/��6k#5�4v�2q
=���l�uo�/L9�b[e�����̯z�ƀG��Є����d�NԸ[��6�Wӧ���{[�L���5�n�1�U6 V�|p�X�⾆���Θ�#������D�#�p�O<����5�E|1~��ͱ+�7�^?�EX/��ǿ�U�-�4-��0�aS3�@��ӧ�+�$�
e�I����U'�U!jqj]2nݭ�m#+�����c�4�Fs���ރ���e�$��^�x9��*UF�韍����Mw35�,U��r$����)-�Y�p#���{�u�K�,t5>�M[����^ԑ�{��a�z��N5���s���x5�q�><��68/��E��F?�oߦ�	�Ur]�}�\�UO_E5X�-Y�f����}Ʌ~���J bo��(��DD�7�뢈m
#3'y�B�J�I�9C��Dr�l�s^�0棹�{U��0�wDzM��� �< ������u����v;旳oߴ��vϖGj��=v_�����NKň���$oϗÐ �ג.���!R7D� C��ex�ǿa�p��z��yfr�*���`k�}V��N������Gtoh���-`���%�N/���4��_��K��/�^.s�耕���%��hu�I�X��nL�u���g�6�R,�>�{԰�.�1�;�4�d�Q�]:�0?��� #u�_�v��m�I/~��DaER]%�A.��υj�O�ֲK�>s�ݛUU������77�Ϥ�uț�?'��<
�j� ���%�G��]���t.��ːܮ�^�fߛu����ԩ]�!��~QI/Ĵ"�ވ;Ʒ�rD��\|G�V����?_V~�w5(���k	���_����c�����������~�ߏ���?�����~�z���F��ܲ��}5����{�	x�?��d<F���"Աd������QgϜ�����=Q7r_'����^k��b@��]Zk3$�m���`PǨ��$��B�4_Y;$��,MS��rjω+{&�"�M$��c/i�y��D�vy���oX��b)>�48b��k꽋Pӂϻz'+8��/���z̎��>\���Q���?�Y,H��@VBM�A�⧭wE��L���O��61�;��sF*<2�\���.��,��#�5N9S{F0#L��O�ч����|�9!���_[(C�;f~o���X��͏.���`���7�@�{~#��M��kpKt�u����Tǵ��Ϩ�*�^��DiE�%y��fGJ�-�6~�&r����=ﱥț��r�����,�y���;�	2��������71	�\hLa�/��&.�>Pݑh_*r��m�M)��k^���"rY�J������-bm\�������hB����\TQ.fJ���ٴ�/]�2�/�_�W��v�\���C{|+��R�H��ZΔ�������zXLaޱj�?<�s���/)��X�}ؓ����	^̮rQf��k	�����}�/<�4�i����_���B7�j�0)�Oo���/A�af4^|����욯ƕ��W�8���Q��U�r�]�{�U���Tj�8W�>�^�]�Z��p�3��?�͸�9vL��#h�-u2�W�
m��l��G�fv�;�\lx�O�o�L�������W��G����n$�F5��qa���W6�J�:��m�ae��t���u�r�� 0�8�t��s�^L��@l��u�u�:��.�&7�z��A��a��/�z����h��܌n�>�!���eei"5��C��[3dQ�`��o/���2�X���g�]�2\���N�;`�5��Sȓ+PL�cT�G{G���2+i��d�`�������?.�W}�f��(�b��r���Ć����.�	�����5r�~�ƭ��T��]#��:u1��Z������+wjB�L��].v)%=�&�C;8�U�e>tG/|e�Qs�rًS�T=\>��Z<�"����/�4j�"���Z��t���S<�%#�D��q�j��>]���Z�A��'�C��%�h���(�����$kQ��� �D���&�~�`��&-]#��\HG���l�[��4��Ы7a�o��m+!�x�Ջ��N�&����4h��Q�"��j�W9_�ӶR;a.�Y��ġnZok��W]nl 
#_��%�fT@SUw{���e���*x�gZ(�f����
f�e��5-��?�I��L䉔5z�����fx�R�KZ����x�)l��5���� 
�WjS{a�_�O���ܛ�;���S{�#�qD͞į�I5oe��r3�֪���8�l�]�cba+���B?XM�'f�vLˉD�0̅[�9�]58/K�ay�E���,�j�U���f@��Q�-?Ř+ze�6��q[�?|��/R5���EC�/��-��� �2� C|JBw=����vls6��$��԰<x�.E`��I	�}`4ou9#�ί��o\�K̼��D��'�m�X���&#��8��C^N~f{�\��Q�,	m�}-ݮ��=��z�T޲��$["�=�r���Z+���y��%��Cͽ�-Z�J��Iz��ݦ�H��%�ư��.�8����e�l9��"sS nQ�i�Bw�h�ё����㱘�_?���P���q�� �o��iZU��rގ��n±`� �o��Py_R�9�'|<��@D�	����O�����r�'�6Pِ��ˌ��n6�ij*7�7lpBȾC�ø?L�:O~�8�r&	Rzb�q};hԝ��bq6E��K����7�f���n���E�4Ʃ�FQVsaL�t�v|�j8=� t�q-3����m�h���N�\�z�\���t���7Y�����6�Ӵ
��@1�NO^�|ޝX����a�Y	�/���] �M���	��w���7��5��6�¿�9��o��7���ݒ�1��uMQ7^��^������/�in�>��>�Z�?�^���0�}P�n������/�����)R����m��k�6����H��<\�� ���x}{E�iL �XP�9ܥ�S�:��w�V>c��BU��7-_��Y�ϧ�ǅ���? y����~�� E�;�6@/Tyf=�?:Tje\��������謊�$��<�Ǭ��������G�Sc??Q�6���?B`�C�D��pg���q2l��.�~��2���%��{h�(4JB��(�{YF����J/S����r��w�@]��z��1]]�\��1g��h�e��Bb��փ�!��?/�v^�6��i�A�[�V����/5�0+o���v������gJ��W�B���N�8+���(S"�s|_0��+W��g����n�z9g⫓�Q�~ʄs��d{MB�-\��B��K�MW<�U�b�Ɓ/a��{�D�h�iQr����b��\�B�\�B$���D1��Q�� N��et_.1���_Hjۮ�3�zq:�]��l�v���xܷ͋(B�r�����,d|�A�T����emw�B#��8��!SGm�U%��R�#�8��)����q[�S�n�-�.��\��[s��ͭb�& �ҍa�5쩢B��1�}�\dzx����������&�·���ޑ���Z���1|͋1��2U�!f��)�����G{"�����DP��;��!�~V�eum|'��4�3�%\���co?;�Z���Y!�;�t p;p������O�!�

3}�P�n����/WU�E�i.(��n� �J�c$��Z��Z,�mw?�A�j�<���r�\�ǂ�NݵP���bx�j��v2�N�*�����0��:����d���@���j��.������󮓍7���Є�>�I{�r�g��q�&��K�}�m㋑0��6�Y]�^^sã�% ���<ئf����!�#P̓]!�%5�d	��B0�bDA�g�E5�=[�۶m����G0A��HO�P��'�O���e@��<��&j\/��#L6Z�h�vt:�#+�o*Y��ǣ�>��ͷ�5]�A����]�75�r5]�#<7>Xδ���	���mkZz�o��&��w�XZV��K�D������8���P��D��ti��RU�d�gM������z��W�d&�)]�N�_�O�"�ޞn�T�*������A���8���]Z3SF+�~�-�p��6S��S��^@�1�w�?�]Z�YPu��3?oR{���'�i�ԏ��m-�:�:���Q�����,����e�J'R]�^���s�"���PI�x`�o�S��	�\�I��eX��)�(y�}��#�Ȧ�Ar���.��$O4�w��"b7\#�����u��G�bXWi3���IQo:�r�c�b��1�84=�H�r�[�#p��e�� ��3�{ŃF�1�]f��� ��KD����Q^+;��9�~��&�U.�W�b�\��0�M�%�z��X�;u���p�惤��MZn�Q�2�ۤ�t���4��!>�pi���vm�MѰ��@�m�okT������y�>&��%�1A[ZA����v��qW�����6ǽ�d�H8s�NT���J6W�+w��1�R�d{:�$9���x�K��/8��ZV��{��Ymz&]'�sk�Lȁ��������t�t`Ya9��1c�<�a�*� ��M�-���sig��Ʒ�Ąw9;��H7�]�=YI���t�E?���J+��׼�r�ϟ,�t1�J�	ty�_ENI��z�x0�Ct>մE�,�P��i�["��xX?I���d�`��6_�������K�������?��1�b;Y_��6�okoh����oQ^�V`����1��e���Ԫ[��]%vXhCy��z�{@�l�ʹNUb���K�p�����oZ�E�Z�f�V�n���+�J)������
6�sl�8�㻣�l&�쉣�!gC���q:��W?��0V5�W������E"7+����
�Cb� ���,�9mR�[���ݲ{�o�7e�^�ͤ�(��d��!_/N�&׬c�&٦��3�*�M&Q�'l������C�w�n�TG��1q��5���DM�y��5f0i�� ׳��1�,���Q�
�_��4�F���~c����\����6>;m�i���6Fo�SC��	I������yե0�`���;��4=���HЀ��9�#1���/!�w=��`{.��n &*�/��U2���Ӱ3ig7b��گXb�bc�����V���%{�cD,8#>	|�(Ӏ��՘r��aʟk���4�n��s���C�Z��1�ˣt��S:zl|t�m���ʵ>�@ڐЦ���M�P�7������{�m�ct���>B�%�ٴ�.g��h� ޔ�ؼl[}����2�0e�O��fw�ϥ����9� cV�E&�>�x�-nߍׅ�h%�
 ��a�ܬ�E/���Maʒcv`yG�-'�`�Lq�̮1yU�<$���&o�(�΅�� ���-��$�%�N%G9'C�`-������Y��.��ECp������8����U�?��nw��d��
�����Jx�C�{B��e6>xTM�/��߾�0�M��p�K�Ʀ���n� o>�ax�~��ݔb����=����<�� ؼQO��=+qs�Yk%hg�R�����l,S�b��o�U�<\����o��S��ȟ��M�-hq�l��ܴLL�R��X�][A���B+<�����Vc��5�,��h۝`#i_T���AGK��Vt��}��{�rtDBR�$;%��衏��� �a�5ϛӼ��j�;��;�abp�A�V���~�������-��	L��Z]%^/Z�\�*��Z�x�~M���y�@��1np���$���0%�5�������]���?'���f�%�7��z�ѳX�o�q�F���I�o@f϶�;�q VU�@��]��nPu_�@\�'WE/&���}�5ƃ�+pL��'�B��2�����r������;���N�a�&6Uq�{�m?�o{uDɳ�|���tzL��苨82+o�v�Baoz�`�@�� u�0���b��W�z��D���U���'"9�w�[ԫ�.Nq���di������d�2[�Nnƽ#,�̲*C1ꃄ�o��;�����0�'�݄��ԝ\`Ru�E7�m�"e#].�{[$�O�eMg�MQ?�Sv;\�j�dP������2�*y]�	Rɍ�Ó�	I�X��"�s?�7����o��F�v]�����y��}���fc?5�<K`�{�
�d�HӁ��e]�&A 1��#=�o	��(���`�3����Y��1�Y
4ܰw�T9_�H��ݍ10\����%vPo.an���D�NƃӍ���I�E��5Ly�!a�
rVL�^�Hvx��J%S�����)RHy�܌�����)q�}�"*�M������j*Y�?^�%�]�v~^� �~��i�P�V9�\�ĜxM�{;[�2Q2�Q�\ @R�^�e�g�U��jƱf�&�M���6nH�-��\�7㹊�$����ʲ��ɦ�b�=.��E�<1j��u}Co�E�X�����@��Et�7
C�4$�����u_�Z�&Z���	ZS�M�^��tQ;�Ά^ÿ��v�X���ޞ񂖋�$�Z3�ܰvv8r����'Ԏ���poJ��H��'.̺Be�����W�~5���>�H��\�d<H������� 8v#�AkH,o���D���#^����o`�O��Z�d�as��ôF5�ީ��.U� �vk`eBF]e�/?���7L9ɯEOQ2��]w�l�zE�%�MQW v�3��4�i�R���d
�e����[�p�|P��0���G��7�}���F;p�ob�ڍ�>%�V���ז��i;�ڇ�ə�%#ҬvH�����(>�v�l�O�f�{Q3��S�X++�� ���([2�����ؔ�Y��)���Z	U��٦�o���\^�p��p`��&���֍�2��:3%�V����Ԥ����!!���ۈ7C�e���F�����X��e8��f1d~핥s�J�i Jd6���(��L�C~�
�N�ץE�4���H���ca�$��8~�qri?�����<̚��1��K9ylh�)�&���h����O�*d�4��Yax�MC�
�mf �q��ݩ�;r��1�Hu���#�"��Q����KY�\�}%�}��.!xt+t�~6���!��-����J���.�Ƴ3�NTA\#�f�7:�����u�J6���8��纜��!����s�&��x?afDd�TFCN�#\ْ|�{���H���|����'jMO�5�Z+1�ؿe�j�Y}e�0nW�U��Ƌ�,�$�|�>�%�>�i#�>y)jn	�&��niN��iDhRX���� G.�����@tġ�G=./EqF��g,��*��ɍ@F/1�?W)/E4y��_C�0��w[��8���9��6�|-~��Z�EOh�*䔏�.�$:3$����C�$l�0[I�E�0�iI��n��Ʈxd'	�"3�k�h��ů�v����CMV���q-3g���	wbz�A|�8aj��KbX��2�=M\!�F�.p��pjA2b�(��FH�� M�~��k��^����%JJ� eС��[�)��5(S�mS�WZJJ�8���(���N4#ޜܾ���K�<��%`����Z+��#������`��3�af�zF�N��֋��q�,�[��H�Į�����bI7䮟FH�	C;���B%�4g����61D�Ǫ�w���clG$1ʼ}����&��\��d<r�A���!,�$$�F��ɷ7�v8X��:�E��ߚ1��U�*�!����]׀&�)�y<ćP2-�i�x('�GQu�F��w&&�0ٲ �t�e�����X,mKI��M�:��������'a���J]��(�8�O�-�+�o�����Z�R�/�`>d^#6;��+�]�|O|n�`��-��Er$��J��.:+������|b񚘿J��H�f�\H���b�r�J��]g���s�7+\ΦJZ�2e�oVR����7����`���c����c��ذP���Bt�n������~��n�C��G�v�N̦2mBp-} �����Ǳ/j � ��nݍ>�J�Ϙ��Q�j�!u_v}������ ���'�סX�)ȵ�M��O�N(>��j��e&�� ��e#+�ݴa�z���g�ŗ�Ѱ7Zg��2]@Ӥ��~���vπ!Dh$�'��3#�J]g���KV�H��ã��;�V^@MW`��3�5��~�	���x+����Ճ���X���(,��!�_����b�r}��Y�mr����d��-�F:�mA�Z�p���$yo���-QӢ~�`a�+?xǟ0 ���9�5P��j���y�a?�H=n x?|3_���rb%���e���`��\�#������G�f�24�$�a�ċᾀ,��pl�Q�j���"�v3�X�	����347��W�}�ي��s[��Ԛ��;�Q�XP�T�����cs{̴y	��:jqѳ5=^�rǁ��u��/w���p�����Ȍ� Pn!Z�7���W�يE�C�bEE�Ǽ�L#G�x��.=5�0�������%�~6먇����F�a9+ݼ>\ݓ���a��@eS�����<�2�Z�����¦cĳ �����q:'0h`���$�^�/ʼ���)��P��+��\��f>��-�*����̜s�H<�����'��`��"��^�S�1N�,"W7�E���`�	��X�2�*L�a�}���F�{�}��ZVe�_u=�
�g,���0�&��=e;��◗�P�H��3|�w��\�%
�bv�`J��^���`�2�A��֚�|�P�Ա:�a�8,
�]R:���&bUab�`]�ƶO�j-�=K1F���GB�qU#<�++E�*`pV��Q�5x�#dĵkq��p[	+�/ʮC%[T�˽QB���R���@�J	�ׇA��;�E	&��j�����6��H*8��Uݳ��<S��e��7��VĶJ-Ω��Aj�@�����5Q�tB�$c^t�@�hA��n�6���+���M��fk��(�H^�5��}C�l��7�� #�8���0rd.'ZF�K"��c$�����Lb��eՄ�E�� [a�k�}�}���z�x�|¤����1{�~���g?`�8���;�u"�> �q�N�0��t^��K���	B(��V�M�pR���I;:�j$9DO� ������xT�%Io��_䰼Z�xz��������)�E� ����\B�|	��" �@ ����7o�(I��g'y��6��m�1�vPe�\)�V��M�*H�Ы��z��^{oY 4�k���>��3��eYab�c9�����N拘���b��q��J:p	���wk�ܨ1D5�kw@��(��91%�z-/��F�Xo��1�>��5���F9�Zk`o�S��+<R�"ho�	?�
7,��Y�ȁ~'u��*r��
h�T����A��������h�+�^|S�D�e�W(�t�Q�0#�`q2�c��dNx�ؾ�x:�U�H��!Xh[ޛ��)r��~�I�`��2ў��
�jE7;�~��2��$o�ްP���f�|�S��w��
� �S���*̓>~���K,��2�&F�k@L�"������6Xc����ɲ`jڙ�G�'��D����ب41"X�6=��G%	ψ��`&��̤���/�"��&��v9�`����}B/� ��yQf"��6�7�����k�yyNs�]��G�n �\Zz�xO�'�yjl���
�'jί��Ѝ�cqF�Bl�;W:�ܛ@����b���F'��A�N�CkBq��8�Qö��0�ʒ�ѭ`ʅv���5|�>=�S$g8�a�&��=��>��S��퇸�1]|��M�X���ؠI��!XV7}���;D-i.qQF����wE��k�M1�oBya��}�
�c�BN�����̏�7��S��ߏ�W���}��V�|�W� CRl�j�V��'7�x�`uI�z��4*�Q����M�Y3�*,��B��Q��`��Լ��4Zz�ۤ�ˉOD��~Gt��eK��4�t�B(����]�o�rl�D�ƫ\M d��4��hg���!�_�@� ��i����G�e�ns��Ԉ�!�r��M*��t%1����;��J�O��J�:����M�w�/u̡�
f�Řo��_Ҟ4a��ꨍ���-��g��%h敿�̬�=��E&9 �� �JX����L��m�s�Kx��=�(��F� ��B2&���9W�ί�Κ�#ƃ7�m�>'3m6P�U�15?��`$_�mP����
��g�-[�"Ttb�t���+�����"C�k�1"��Y~_�'q�丶�7����F�<uv"5F�{HMx\�/u?_�l{�8��dXUk$��KG4w�q���j_@�/n������G���炣��w>�7�1����ݐ��V�jK�ܒ��Dy��sa��^em=eI��R����!�=+����+XV��췚[��q��l[h�4�䫊,�M*�o�[e�����{�ݟ'��Ow�GPuE�-%�)�,̝��EN�̰A;?���xJ�F�\qt����ϚL �J����o��a�NG�-a��c;�6�ǻ1������-�,�뺁1�F��g����^sK,}��t����n�H)��K�����e�a-?��0P�|�d�N{ؗ��"fv�X;x'���Ό�9α_��Zv#[8�{�K��l��}�Q5�(����t*�N�#�a>3e��e�ߙ�64;6��K��Ʊﮊy�D?�Y1=��3�4�V df6�0}f�7g�Ydۛ7=<���h���a���w�:�S�B�@��p�l��q���&����*����h�����q����)��������6��(%²V2(r�8.SxЂ��4z?o�Y��p}�`E�Κ�����S����h�^��ͳ��3f:�\��BG{:�U*��{����_9ƍ�b�f�P��
ռ�`�D��ݿC��U����B���K�b�Z~Rq25��7���zF�C/d�sU|y�Iք+PHD@���f&��ۯ_�ꚒEǰ��4�?X�{z&L���1�ì0/�y��T+��;����j�KD@�څ����X
�fz��J�n)�~���=�YhG6!�(�d��]z8kz�x��.s�����.-� y�X��t�L���,���D*ϴ}�x)#4,u��(�TyQ���x��q���7����ǕE���uVNuN�X������Co��- #��#���#? �A��q�eH���Z����Z�P8aέ����2�NAs�_�j�_g;xK_���{��/����/c�ª�ݠ/5;�2X�����tߡ;�|)�N���w�S
oJwD4:�rTfN|�E��5B�WT�<ؙ������X'���ΓE��n�
i��k��#��Æ"zsw]����/�<�s� ����([����f�p�ه&g/�ȇ�A[E1�>w�[8p�}�l���3N-"y�t'߅��_��x�ܨ���M�e�i�����8�E����j��%u<�ͻ_��?���L�k�С���;�J�6/���0^����7�'~s�a��v�~x�O֤�[�GV�e�7g�^�ΛG����MᎰ��Ǆ߬�����U�%����W��o7���Pp��'w'�d�j����o%3���dl��+�3����vr�D'��Q�{��)׎q&��H|�t�7�I�.�dw���RvQmyd�p~���s_Ů���w�s�t�����]s����v�
�=�B�!St��Š��?뙴���z����i�u��d�lNM �-���T:�x��-�yBc󏞚�ޯeT=�VWUUj��?ک�5��3'f����9o�@�!�_v<4���n뜥I��g�5��B<��^l�J���j�gP*�J��^�5�!N	"���u�Ӝ����������z�w�1��e��n�E1|)�U})o�s���qZ�l4شR���d��~�/�0X��,�D�i�u��F�]�Q��F�#�YĜ�%�&�����P��O홟�����t�wt޻�f
�Ea�ofEv������T��%�c���:{���Έ8ģ[����ךª��J��rL�+�N���Z
\ԉ@�F��}��)k;b�t����wz�.�4$?)��<��ɻ����w
o>�jѹ)=&m�1�S4m��~�%@:AD,˫dc�����Zz��-��^f
�I�d�����FX�YS/!H���;eg��Ɨ���Kۃ�~B�P|݌o�2�_�lKCy���s����]��X�Z�W�����C:�t���҃�d0�
�b�.N�=�I��fzk���5��\�B4��r�8s�e,�$^����l;wYTHPtX8�CE���e����,�6n*8}뉟G�tJS�0��]�[1|T��YOu��f`�˗e
="w�e]�w_�B��5�|�v�Ts!����F����">x7��dP���PG��4�6��4+�69�'{M�s9g����݂�a���ԂN����t9-�|S��L&����ҁ��j����3�O��q�����r�)kl������-�]��J,����ٱO�I���{��p�	�$u7X�:���
�W>��m����m�"��Q���ck�a9�V��Y 6Yl�s��=~�b�a�oS}�yƪ�ƌw�Y����NU�0��5�
Pex�S�C�i��G$�����;eş2ݓW�c&���.�6k��I����s�%��z���zs��X�"�Dq�:\��(���a���3�\��0�,�:V��p7�XK�_�<��U���F"��mb�T�tT���>1>�^%*����Z0R-��a�$ �'Zn��ʏ�0c��~����uq����tܤӄ$�n�Ġ#4�oYN��H��.Ȋm!|8`��l����փB���s��'�k�5p�D1=�f����cNn����|^��G�/W�̌��r��Bu�����]'_��DjE�wH��?bg�J�%GǬ-����D#/�]�oq�hֆ��,Hƚ���՞.i���4r *R;�����.�0\�������C��˨ҋ�8�Ӱ���ؓ��3&(�ƣH*q?٦��;K�	-+v���0�~��Ȅ2���=�M�2RlB�k_���cU�mv ���h��x8��w?��"O_��6��!�[�J��Ϻ�*���O%.R}{xZO ��P�Ns�؎6�֦j��+�(����bM`Oy���>ۈ��p�����:}��|{��o�{��s�a՗�e��@���Q8֕�؝-p��%�-��46��yd�� *%��ĝF �r���=�Φp�$� �.���nХTuw$Q�uAa)ɬ�"9B���v#>�a6�ch/�)�б�#4k�nˆ�g;7 gx0��L�P�V �Ca-��G]e���>�Vy�:�p���@kP���~�,9|d8k�v�q��9����]�n���g3xdi{B�k�v�q�<�N��/D�G��߾�ΣP��Z���d�Q��$�s�b��w����@�ԇ�M����IdD�����tjR�aS�߸��>��$Z��e܃�f���e&V�#��$6\3XB����$�|����SWD!?5&f�Tġ�����	~?r�`Z:$��`k��9���h�N�,m�������L[�����1�sJ����xG���+l*�$Ԙ8L4�D4�9�"B�jj�-ְe���H�Ь���h�uL���K���Q���׎&~Ca"-%BWδ����}�շi;V������?�h����5擓G�y2�Ө��zDO�Df���k�o>l�����fs��_��a�v������� ��vRf�u:�oº��������nEJn����;�0��&c}i�{��놞�\�}�'1��������F���DFᱥ��}�"r"!L�N�o�S8����b�Vj,�z��A�+*�
�/�ɳ9��.:��$��Ȣz���G**  ����K;���Byr�ۋ�� �Z�ϕ]c�6�y������N��� $t�wV�=f�Iė�h}[*���\t�2�禙+7�A]Y�5l��M�onZE�#� �G�9'cC�
�j�3��!%`<��`C�dJ�4x�gv��/C���u��)"��/A#%wOZwy٧(�i4�bY��-?!�٪���ic/(���$�vP�N��h���If��i75%@���	0%ċ�z���1,@]�t���E:pk��%:��^w�z|�d\s�X����]8�7���z:� ��2&e�V7q���q��o�;㚱�1�<�@�b�TTۏd��&<���G��4�
����(%�`[�6c]s�}H��ج�̮ϕ9�d_�s _/�)��Z`�ۇg���(�����$/	 �w�5R��4E���J�D����{����3�<�����(��(�/.�2�cU��,U+Ԉ��p�l�%�"̍*�H<�;��o��mhFKF/qƵ[��4;�0���˨��ɞ�Uz��`>ߴ#h �����'݂����0���ml?V�"cd&��d���w9ixeD@ w*sAn���6�Hr��Kf�kJ%ώcHHHp~�8��/"qԗ��I4�To*���=�y�X#�����O���)���ď&���S�f�Pg��LV�3�(��?h%Rm̍��>��f>j���t��:�w������S͂@��:����'���0�e��PM�B�b�D�݈�2�i�����t��M�NW|�l�c)kQ|hBΰj=�s�`��<w�X�C|}�h��̂4�5J߇7J+:,�q�vPp\�o3h��ό���D�rN�jUp��3HT���"X�S�j�����:�;N]��V2D�b��@��>�)�8Zo����D�M�8θ�҉r��2rz��<�ޤQo�⒕�]����kc2��&e�F�0�،g3�A�5nޣC�$8;���ѻ��-u �c��hE7HعW��������n�c��h�����dϣ�̍����nc!�8��S1�O�.���P��ZP�� �X �$1���8�a���Uq;lO]׺�r�[#����DS�Rt��,�7�Q&p���mbU�8{>���İ�r�L�%�A8�S�����{��@�5�e�x z9���B�j��>{s\y� ���
ehYӨ��O+�̳UM�����m@�Ҋғ�ŕx�j�}<j��myHz�o6}�_�YI����O�F���W���'{� ө�M�o:�8��J�LY�[�B�y/8�XU�����%��g!�q�o��3��U��?5��z	܏��R+&���_����~�ű.��o'A����%�����PD۽A�(��`�|��Q"*���+��;�&cq/;�4��P��I�A
�bm3�T"(�'��s���'^X�~�M5n������x��8s��]4_$0���0��r6��?F���D2f��LyXG���凌��	�0��$&8L�2�VM�UF� ȉ��Q�)�.����Wdզ��҅T����"���R��l�Ȩ���b�pw��נ�6��I-��94̴j:��x��'��`�Q��PQM��xCɆ�
��d��-��+��J��4P�>����=s:J���o��ݦ�$K���c�2w~� K�=8`�~޳;6vW��))��U�<�vxdmd!��ϟ��z!�BA�H��&� %�y�� �%�
O]i�'2���>aq��@�h@~[�7��=P���h��83��֏��KF��՗	�a�`�S�xqi�F׹���V5D��)���NI/���vQj��/2X��7��Qz����y��#���X�p��T%���>�
P�i׺m��C�ޖ�t~��m Td�ƴyP����X���,l�����)�T�+m',k#A���::VR|m1ʁ/�77ȶBW^�Ԫ'iO&d�G�H�aA�}�S&�}p�2,�g���԰{���z�Ȩ"��tZQQ�*��[��E(��8�dC�Hܕ���,�[���n�<�eNR�hR�4���ݲ̑�7aОͶ&�4a�󬑺 ��1Q����k}�k�-�����6��ZUI�U~�?�_�7���vGjj�t�'쬹�IɎ!`�'_�VҊ�CH�w0o��M�s��J���i�g������$Exq��k�ϧK�����ά9�Q�0IKN�������K�3%�;p���b�(�E%Y�](��`�)W�O�K�O0Q�s����>@r�0	�ҚC7�3$�Z���e�*�����
�Xj��_Un6�J1�!�^6�Q��%3��Ib��<>bg��W�PmD����@��<��VN�7Z����M�	�"a#��q��q��Y�rm�Q7��$�IB��$� �ի�9SV�J���$�%W�&�¥i靉%��`�A�&$9EfI�@Q���葬�*�;�mJ
�9�_���K�W����`Z3�&��sw���]7�Vj��*]����"�1�	0��������T4�c�����j��x�[¸�\�������̽ H:��VV���$�_>$<
߅�_I�k|���N�T>73e��fw#s��	=a���mg��ӗN�u��.�2��Y��*���Z��KT��]�E�;d}ҿJӜ�L��#�ђ�Tn���|'��r4�`)�ST)O�ϳ��=���aq�;��
R��9�B��$^��W����H-h[�rZ
�s�O>����t�Ǵ�4O_T�^UF\��25�0K��#V�fB� ��'bl��g���]ͷg���_Q������'��Wi�B��fӧ/$*�v?Qz��~��g��z�W�%��J�3����W�꺅��l���W�D XbZ���q�_�y�D�}_��Fr�W��<V'�h0��$�`��5��2�k�UQO����Z걜)�[A��InmiB�A���gmP�-v}��E�>�=ߜh��Ј2�&�DJ��2�Z���o���a}��4a��8�B �x2f���
'��Ka�+���Ԗ|cGɇ���pZ�g8#��U��-����,�۝|����x<��}�c���rY��x^��>Դ��gW�໋��\n�����{�qXdhc]�+�.�3��g{G[0ؓ�.&�})6��[ԫD�ڿ6 ${�G��&$E&9�y���:���۩�?��t]�gz�� u�H���Ģ~F�\L��t���c��ү��z�����c"V�3��v������K%ݹ��y����՛�	nI��Z�̯+�n�~�F��vY�b�_~]kvM��v�?lw��y%Xy�h�$�+�/���}�du��	��˱O��7�	���>E^i �<`��4�o�O�Ǟa�\�/E2�]_�q��.�`�#4�&�~��u۞o��~;��42����ӕ��lNl�6��*�nC��y���|�>]����O�]���G�
C7��\�з���T.C|G|���W���W3�/ë˿�H�_��YtϿ���5�Z�z[-�y�Q�F��c��p\�}����2�(l��[f�O?�*��kzu��(�ԇ%biJf��i����?�欎�sLg�b��r�Hk�4F�*&=�~S���U�fڒ����W��7}*5wK?�$��6�"�x�>7I_���}Â>i��j�H���zm��6����t�����O��9|)�m?�B�u��fٌ�^�Hq=����P��`��Tg/��6�
��Q�:����q�z�O�Kq��%_����:w���m�
�L�L&��<��'f��Zr�#����߸�}�R�Mʃ<�)�Y[љy�f=���E�"�b|������l��Jz.�t�k�m�����F�X�YgR�i�f�_�(;�����/+��j�O��H�:Z�`�i�>����l3'���O�p�r��x1���듺Vľӭ���W.�l��N���<�T_�ebſ�%�Kݪ�ӟ�:?[�����y���q���o4��#��;:�]%�v͙������s�WKN^������{�3i�_�i�G��ŏ��B�+.���C�\ѽ��{��������"U��Q��?����*�0y�jox���mi�s�zi���[(m�q7Ι?�ྜ�/]�����n,'��c&]+���*��w�2�&.�����.p���܀����I����_����@7���܍d�����
� k$ʴ����/ٿ��<�~�ߊ��;�b��q�(�7{����i��*�RP����DJ|�@6�ܮŶ��bui))���S��;��^��p�x�&M�Ih�p�n��.��]�c�����������->��=<�����{�֢0Ԯ����wx�+�_r�9�5�x�>��ޖ�
x�N��HoO�it��4��s����;,�ly�W	�	wa I����r$H�(��.@�р�a %��(��h G�$��9M�����y�}�N��ު:���:@T�*usO�~�ѵ�,�?��*;�*[x �o�� T6�0Pí� ��������;U��ZÜ�[�,��:��׉.��G�C���Do��Q�G�����R��q�tt� x�;�Pb���\F�B�L��s�;� ��]o^����|�d�c�L���g��'L���� 	 ��:o�^�3넞�����yUN	�Yy�� hE���ĺ|}�ɺ�;3H�roqۅ��bA�)c�yt�.-N;�P�U��[G��kfg��r�ׯ~N'ܡ�����
(�q`��K�2�':��=���p'@��+Z�)f9��Cu$�aQ������?9;=lIa��� ����{RӜ�3)���!����ˬ��"��9)֑�}��I�2Ȇf̭Q)��S�e���[�2+g�W�r�����n|/���v������_��x;�[A�����2dnb�<�a*�<G*`���Э|�F��L
���Tj$�)1����S_�����c7қ���aD�f���]�U�면țh�	���r،�
�����@9b�=2~�4D��j�Qvc!^��N��7�-fh�@5��l��.�b�ܺwRA6�獼-����|Cq��V�e���֒����$1� ��h��w�H��)�%�@�^B(4����k����;�7��"��DK�7��Á���*;~�#.�7����������s[�:Ve�Pn��F~�cH�����
>2�H�n 
��|����ϭ�pS�+���:�Jd��;3}�.M�� }�!q� N�6���w�*�;-_x��{Z���1����gЧۍ�i(�cZ��mc�;M���3�o��ꙋWu%a�g'8?֬y�\{~��lJ�Qi��	�(�/�=N�q��J�/�\�����Y�$�{���<O�Y�*�����.A;��Ytz���9�Kq������o'�����A���sO�$�[O�b���m`���?hTO���P/�S��[����[�ͪJA�*?�rP��T�'5���NtD����w����?�L��e�b+�<��V��дqr	&��r#�C0��3��i�6k����6�ͭ���Ke��.\H�jy;Y	��&p�G�}r�JjB��{����I	�������(V2��A��k�n�s�9��V>��M��ʴ���Iھ�Fa�;��	��6�i�Ň�1����5p�����z��ey�\@��M��q-J�y(�F��c���^a7Z���g��\�ŷl�w>z^�vr(�I0d6=->g�P���n�At.dSұ�GW��=�A̒���U�t��v2ׂb�o�0���?M
�mT��r���~�R�>�!��I+������j�ZY.Vw�Z�h`.��JS۹	�����+�s��]��t+痂Ÿ����\���#%39s0W���}����� G� eٌɱS��
6 D�ӽ?��C�F�tlb�.%B�E���jP��a-��
`����v��v��wʤ\r��/+���R؋��.΍5��c���c�|5�5;�6��K�� �{���!`b8�A��	ŗqc�W�!��3���O+��$Y��o�,~j�a��d�	�'��悩�t�nČ�~�Hu\c�;8��79� ��xU͸�&�g�Ip�I�Ӕ�Hv���m���4�Od�����Y&%�D4�U�*�h��h��z��<��c�hDX ��4.z��(��&�9���$���N_?�� �<kg�_�v�u4��h��r����\��u(d�2{�����;�ݭ� %�ƋAs��;��*�L2�~�5�r2���B��S;�}��0��<�yğ5�z�i��%�)Y.�s�Lh�PxN��8.��_�`�A
i�ދ�����X���o߄Mas��������L�[ɠE�wD�"��5��;x%��v�k`.�d��<�F��"q���2�V�S)��}`F��� �}��:�T����e�-��s>�Y|�̷��`=�Y�7.�6�} Ngf���0M��t�w�t0X��&�ϾZ)�"Ϛ/R�R�z:ő&���-1�Á��r�F��[-�o%���+��ߠ�`s4[������7Szۼ6��љU��Q���+�C�D"�N�Z�h������f(18m���:[��?�<�j.� ec����|P�(a�(���J
(��	��tC�3�[���6S��m3+�ZB��	�A�/Ո���*�#U�-:2l�-���g�qb��C�
tR��E�҄僁�ABU|Z│��i�b�D�����m�+ Y���.}RJ�x>����z�����Rb�4DI�F���?��l��:���`��y�6������8�����7��.�iWwق����ގ޸�K|����ދP��f� ��	Ɉg�K	��F�N�����FU�dYQ�q ��0��?�ѐ�q���<��r�CY3�K#v��S�6(�k2��&���:��F����o��s:ڡ�[a����m�;��rPUJ�mZ2�����m*��.�g>�y���9���dV�թ�����F���kxd.𐝯��G��o�V�7���H����z��="m�W���O��Ok�t��1`��Xs�6T{� �[�X�}]��t��F�s-"��DZ[��8i�>��q�nn|�;(�i!�5�r�n|�ج�TX^�6\��]<��(~U��%��c���LR�Y��MU���ٗ��5zv"z��?ƪڃ�� �~����һ\7�i%��'Ui'���m�iH�:�g)�����Y���7�# ������=�U��ϋ͝$\�^���ެx�گ���"�ZQ��bk�>�r�����@��6���!��3�iÊs�X(RRU��^|�"�=���!we�9�v������t.�xk��bk�Q�z�*?���"�Z��¢*|lE|ޓ_���ά��|���_��QJ�yJ�:׭MM��,�в���"��t�� �n��(i���֋j�b�CA��,I���Vy�A��|i�ib-	��KF>;)w.��ֶ�&��H�4?sۛ�$�Ȩ�����~�wP��?�N)���S�Tbŀ*���e�=g�&LISp�CQ 'ը���j�6��~���/[�������X�=���.q̅�$�>�����ԥ��
vw]����0_�+M:�$���x�t�g)-��c���Z\�1m�[ރ\9�
�h����7����Ag��r��mΨ+}�Y�s��J���Ѥ�	��8L�f�5�a�Y@����ǅ;���hc>Ș22-Ͱ�Z�9�b�u+f<��8 �|#��
[��-�{�h�z�ɒ{��o
�Q����`�V����?y�ކC�v�9?��&� ���p��
�i�7	m\�Ǒ<8���#t���<y�`u�I������8�(����Ҵe?���Y�譣,�)q�C�Zc��"��W����Z�A�A�E���a�K:S��CBd���	�Yo��w4�F��8	���|A���#o�wc�ޡ"��� 4���}JQ�������W|�Z�I���`�^/������za��k(��<][U?H�:�5`��K��������C@b�AZ�˰Lǭ�#�?�:+>pNj�?.��������S����-��f�99��aNK������Jb]��@J���y���\ ��[�a�ʣJGA^�Np3�G
oZ�#��/�3�,��XcF}�Tӕ�z
t�u�_O��Om������p�W;�O���Cd;SR8�[�~Y6BW
AZ-����5���iJ�M����h�����[|&.[��}���Ե+)E���{uh���4��MVJq�W,W�l�x=w���/���F�j�E���+�HH�QT�9`un\��{9Zcjm�]W ��ӗ0sQ5�-97�,
 F�k�l\��=U�"&P�'@�_��8郌���2�䐌x�|�6c6���ˁ�����{�KS	qQ�����t��('�T^P0�°S.T��&"h�55>ϡ˴�Ѳ��j��j+�|��P'WQ��.��O97��V��B �W ��_��/rU�G��2���3�,ɝY������
��)�bNtf�m���\�b��;Ԭ�IU q 4�di��񦣮�����Pv����EF�Y���ncb���څ�=]��0��]������FTN&���>�+�c��7r�TӾc�R�I÷�⛔o��͡�w��0��56��Mb[��i�o��,�$�3kȟY�^��[D뙔��=��ː֩�<�)6*���q��7�f7㮕��X�NxZ�}��������I��[S��+<3�z���La�x��&�wy촻�V�K|�!)����A�A�FQп�}�u	���V�y&��� AbS�y`���$���z� �P{����ܛ�O�C`�G�IW^Ć����C�E����V
�Ӻa��$�&���Ȳ�~%� z@,������(��G�z�I�S[Y&��.w�7�$���~�jY�=���t��h �EP|�g�6�5
C�#�B�g۾?12}����K �*b��9�����]:�ty��"��{�W�l�\b.�l��Z/�Y5��Ż"jf.w�����C'���靕h���)��蝄�Ût�+�z�D;�(��˛�j�X���Ȝ���c���
��|Q�t.�/���]����9
��I��lX$p#��l��:�f���*ķ�0���\�ֶ1����xT���c�t��(����Ǒ�_6����JUwz"U�g�ޞ"�r<B:*���b�Ý~�7V�)]U����ƏF��#X�b&&-`Z�Š�����克�p�2[���j�����`�LrMԲ��+/O6'���t�.9�A�] ����2Uv>���n;���XI�h[E�_7<��	���$̣T~	PF��"�Pv�� @�C#���-��l�A>�`m4b|��I��T�ZBKH���E��<s�pʷ�+�uLfg
�hz}�G�5C1�Cn��9?���N�m���$�n���ST<�̍j�!ΗsR�����H�t� ��Xnsb�{��BPyԾ��le�;�0H���p�g�T���>te �.TauδxFR��gq��X��b|N���**e捊����E�b��4F]:Ɨ7�tk�Q����r>��Ƕ�'B� %:��_M�Y,=���+�yWE�j�m5��<B(��K{��	u�2���Cb�<�QJ`�M  l��e����x��.��m���K)��˭a�F���}ݵ?�}g߽������'��ӊ�K�f����/�"�A��V�����ZϬ|��y3�T9�;Q[WY�v��V[P��Q�9}�?��tc-���I�jhlUFWڱ�|��GWP �turZ�b�+@e�����#�tn%��Q0�H$�#W�n��O�MhBH@��a�]"�ߒ���L2��㝏2�އ�VqS��1�EaŘ�SA�][�Fy�|$����B�h�Y�a��� �qk�q�ڣV�w���g�@�s�ܪ��3�N�~��4�	�k`e&�j���y�%P��
�r�e��u	����%�ǩM'T���ŌV���xz�ʅ5�L�*��ހ�tCVG�t3O��N��ZOb1Te�k5&�3����G���of��`<i �-.�9�mk�B�r ����
�U$��?8��ip�"���N��R�*V�ھ5�k���wS6>�-�k����3Qk\s4Y�/�a[W��1z��M�
w�.�{[��>�<�L���9��Z�G>{�������̇�&��Ε��߅� $��Kj6z��x�LT�,vd�nG��T�弾�-���O�k��.�n}PA�-Y��{;�V
�[xԡЎj�ۿ�(�݊ �]^���Ox�Z�44#�ё��Trb%̟�ڣ���?�k��k�+���T�;���F/	-���o�kY)w�z[^Q��HS|o����|E=j � �2(Ot�la�X�*�Q�K�!*�+���ՊX	pʢ
_ N^�9$=1O�`��l����tZ�U(Z���a��)�<}��z�ud�34FK�f�Ǜ�:��͍�`��x:B1w��Mq�K�mm����V ���<�2�?%����\�����<Z���#��'%�A��5P�o������/�BW���p���9����c)��A���咼D��皩Ϗ:ax�F����2_����3��I4�yi�rP��OpblW��/�p�|�(E��1�`�S�Nv'�g�EZ)��j2޼
�%@��sR�*��6�j��)t�A�h���;��f� Qy�N��z�i<'ds$���8������p4�hi܉ M��[RC���(�!�G��<��zƢ+m.�×�MN3�������z��Z�:��)/�GL8׺��\��{��m_j��c
�]3�S�}M@#��M�oޙn����~5AO�Qs����[j54eՕ#��+M�x���Dᕝz�|(�����Ö籧��
����}�����
j_.�_����WS�b��6ɵ���g��Q�E��΂MT	�]z`�@�>���F��#L&��BBg�V�P�׀TF-ע�/ݶ^xE���&j���~�����z"Tw������ m�x,��<���agN}k'�s~I�kc����2tŭ$���<,@�^4X��gsm��ڴ���6ir2Ci(�cy�]Y=���4,59M�s!M&�u�j��į�"e�˒��E�s�y3z��[g����JW�f�<�$Ԋ�P�O"����i �g�����d7�=G@�3�S��8-*��nQ㓔��j���H.���E�'cs�a�1��z�	%��:N�@7|����S���qP)2"N	۰��'���T+���D��P�W������j�!���V�#m��P��.i���Y����)����]�e����2'/�2QX���uTr�^�B_���l���|CGZ�o���(���9�t��4ڌ��KkA�0�\:��J�5�[����(�2�R��g�����k��we)OH̉Z�eT5n�V����\���܀����&�5�`y ����k�� ���/uG�l_�$޿ڙt؄}#tk��3�JFX�/�������Hxx83���&��,��9�"@c��đ�#�QCPT@��ϋO
���[@S�����g��r�
�:M���_Vv�* �q-U�hk��U���}U�����:�*����'��JrkG�),����p���OPHXC�� ��?��?�&>d<+}Ғ��,�r�}N����������$hz(��d�8�a��p9����3;4j{�l�N؄N�� "��[���n�6`�nV�����uq�k�����I�j�ZOc^Г+z�y�=w�خ�63/>�DN~@*���0��
�b>�:��i����/#o�yJ�ƻ���X�R
s�)�}a��Wl�?o��ZF��7=��E����T���
��!���ܾ̩���;~��<Q Ϭ�������B���cdq3f#_��yt�q-�A�3�[�� &�@,���Е��釾���<+�4�0F��ǤrZ׉'j{�|�6˖Nz3��;Y�ؤ�6���~�x�*<+1�>kW}�x���� ��;��* �QZ��!�
�ퟎAVg�}?�_�3}��}�o�k,k�����:���<�6�|y���^�D�G���i!zWv:����}Igޥ��޻��߻Ln�;V%�AW6M�=P�T��e1o�r�t�H�0���F˩��8�ƞ���}e���l�es`�����N4~"��~D3�p����i�r����Wֻe I;ɛ#�?�3h���`��B�<��xG靾�Y��i��S���t������������Ç��#��on\۸=ul�
���V�^yn�Υ��N�E�<�jN(}�����Z��|#�Iۉ��G�d�`P�|ƣKf��&&��m,E9 ���q�s�i�OB���})�f����ܓ�Y��¦~� �L���=kZdk��I̾E"p)�G&Eg�/u�Dr�r��o�2~�$���k�SY�,�X?��s<�����T�:�S9����~hzϖ��/t�2T�0��H0)�r<`���BT7���΄-J~h/���|Z��)X:��)� F~s��Q?� �j�E��pg�>\V������f�$�-"�AWj��ܒg{�5:!�굺CS����@�k�B{}���ͧ��uh]Do����;��	���[�k��꺱����,3O�U�y���Qh��p�"��bOvl@4��U�����^+MܾS���`8��L�NeI��D�&~!�ɺ"�_05��GcC���/�L��&J�~�����-?�S�o>���8|��] ������k+N��w0�׷�g��j�f�90(�:�0��T�Iқ�}:�lP���B4�_�wh�g�����Xv��� �Sw�8P���ߴ���}�����H�L�\)�O�Õ%���?��-�,���LH����ɥ��?h>��KxWc=���-����|�h�����c�z��X��W'�C��G\�!)kwFg4ɻ-є�,��-KQ�o��$�ۺd����{�`�όv����ȃ(1h��ӿ�"(&�7$����YH��=	�&�Z�k{Km=�ki�A�I�nY�y'gﲵ��P�.Y:�r�(C73�2V�(��Y��6Ֆ���M�) @BC�l�fySO����R��L�
w\�P�x���j>�ܫ�� �Su��*�/��ˡ�|�ȧx:��_�v��������g �}?��$*̽���df�&�p�fk���1.���ߡ��g���e.��-�'�F�e��xa�U G�&��{��e�Y��#O�F�����+?��l�x�ч�P|�O[~iWmj�d1�X
����:d��Y�W��#0�����u��}��������j�xZZ���a��LL���x�����/o�5� �N��sa#��濥} ���b;iM��2Y|�j�h9��ՠ�;�v7����9���F�ŋ�FP�ňM�"�X`��J�v��eh���E���2N��oޞ���|���l5�s�e̾�9�N�>~l����{�Sq��ktT�ڲ]�O�_�-uXw@Eҝ�n{'�
�;A�����sE�V
�ei0i��*��1䶢�cxM����E�x�* q���l"��Sϒ6�!�v~�d�\kҗ��F�Y@;L�.�����\"k獊�����o͕@�����]aVi��Ȱ%}P�:��v��#s�ҵ���%�{So;D�I:���W�b�M�
�@��� o� (��STF�s�#U/㺸g�6��n�B�}>a�����tF�Ү���"law6��Z���q �t�m���D0C�^�� �	��Լc= VF�D'c���?:b�ݓ�FU���8}H �;A'�	c��1|t 5VȔ�d��:�j� MTj�u*�qu��V�z�5sU%Ū�>�f�`����-g��\1T�F��K����{Yk˦E3y���@��V�V^XE�̓xw��ؠo����qH�"�����1�X#��Bȕ���?'��,%'&�,�e�S �MN��S�5�B2��Y$[��ϱ����������fpʿ��v�~��� ����h2UV���z��UQ�u#Y�k5��4yи �U�վ�8�R|U1� R�իrn�3v��qq��#���Q)+<�P�O�Ԡl@��׊��$X����}�
�*�X�J�+��;7�!�W��r����|��?wd�:��XB���X=� �Y��׵��EUW�NQ���\TX{`���ʺ��3*���v��j-_�Y�^���՘�|���e�<=�$�x��F�O7�͎'��:}�kE� �Ӭ�J�_�+�G����>���@�V;��� ��	e�k���PD��}�{�`K�%Co���N�=�YZ���E/��PJ���3�S���D�DF*|� �ל�u�����At������pb�u�T�s Fݲ�T���躴t�z��R�P���o:�����`�i�Ykؓ�S���x�L�����Z�2�f7J+��i�#S䷎�&��ǃ{ZP�L� ��$=��S���J�wc��{,�N�D]I����n�p��Ϋ���m<Vf��/^4��C<$�NR����i2b��J�� ��[J*��l�@���@�S����f)�ߒ�H.T��j: �f۾:�g���U�|e����:��瞾���e�%���ST��ݞ>�ڝ��?���y�ם��;a��������_�P3]?4T �8����OvC��R%�yr����U���x*�<�������!�,����m�,ѓ����d�[��.k5��J�/$�]��Ld|Ʋ���F! #	�����.�rφ��"�ӕsd㻟�j�k�N��tg�j�=M{�kS�޻���"�R��.�;'F�Ā�t�1VUKƥe��k�� `��W���0i��b$�nYZ��_���{ s�=�Ǿ�E�d�/�4��V=� �35��Rx����e�EȈ��(ŗަJS?f����~������_� .̛\�j���#d�t=�t@"���dO|TC�T]�b�"Kg�5��ŏ{4c�p���mb�;0Y�n҇v��JS+5�Ӽ�>k	���@���V)�� Y�c�'�Fl�I�S��07��1;�!#���~�'����FxB2�~��|~�����/�#	o��н@ad;�7K���?$��3�������;ܾ۠ ����a̾�F��P6�}�v�&
�7�mZ^ϻ�I��H�'!�3��S�O����gR`���E�9�?�A�"4�O��Gn������2LGC�5�n� ����fw���2�Q��"r.����Y�x��rVCr��(v1��&��H3°'�~�-�g;r��8�_ȕ���ڸ�Y�G�����bc�ul6S��l�:�h���~b���Ъ� )_v,��s4�S�� ���(G[IP%�|R�H��W���C+��f �Z��݋}t��!P���ꇹ�����x��@�˚�d{��z>�Ĵ����T�9�VL�Xp��+3�~����L�F����0�~l�G���� $��:��5��[�ڙ��%��>�1�ꜯ\x�hp�8u�F���R�1��͘�Ud�r
����𤃊R��s��ks0��%�6���p�L����d��CNU$��ڙiT�P������)�k�ݫ�ɖg'��8
	9��Sm�3�Ͻ&�+h�rL~�T�W�M���/�c�A12�%�!�U�s~��Nߢ�u,��"�>�Ƅ�h��ߖ۔�I`�؀��[�q�����Dm�r,��g�� @��W]*+�s;�����/�9ܲ��qI��k?{���A('I��u�_~[>�n��jP�}d��KP�62����8I�'Ȓņ�lɛ���y�AH�;ߜ1������F9��N�\������P���^7�}��-�p����4�jD�zM�A��A���|��c��d��U�C2c�4�CU3�y˵���.I��Ԇ	aJys��~�ct�F�R%�]&����)���Zo�5Kn�������L��z���3���מ�'�M\_&�.z\��)��%siÕNUc�d#�yS�Ut/E �ۗ�k�d�%��@4��X�i=��$�x��8E�*�$�ק���T�춄r*H&�v���l�&�?���Y���?��ťC��7�:Y�W�b��S�=��7�AO
�z�ZMƋj�����wܝE��1ݤӏ���\�ƾ�'GEJ���^��?�2���c`{P��ŧk�mh\�*�����1���ϛϜp-��_/���a�e�{7�5dc:dF
��&JiL�>�+<F`�|�F�;^�5Ӱ�a�!m����0�%h]�B9�Y|��w�TY2�27����"���Vf;���,��ǡ�f0��luhۍ�kXǀ�j&_��CC������g���E���$�8��KM��;6E��Ӏg�C��p1Z!�l��]���4�~.@����~�4�	�%�3}�h��aas���Ճq�u�x�U�6�N5q)��������,'N�rAG�=3�}K�ouQ���ں�0������n�v��+��h(8�+3�i�cjv�_��mȭ���LhL�6}��Nl��me��A�H������
Ŧ�]��­2ܪ��3Aˆ^�%����n<��F
�6w��F9�;Ц�����!�z����x�t�:�=G&>�,N������o�L��w�%��OAx��S�+�/��a���x	^7��t(W�k�_N`[<{���.w�ѥ��0�'�kᆬ�>Կ�'��z1�g��C= Pc��s��^���6GT�C���緖�۶&�v2�-%T6��y{A#^p���� �.��GU3�=��z��%l�Y�6[�h�f|�}׌i�B�^q�����,}�yB��G�mi�D��"����3\��><.�(-

)}mkn�]WD+��;6v�C�=�C���G�t:��& �ڝQ�`�����bgP)�_$.�n�-�;�ۗ�?��g�`g-�ץ���չ�\�{�Yit�a�Rn\ PX��9v�M��W.p`��-�2��C��a|m����2�*8P��,��N��s5�Y�Y��4��G헻 	OgI�T�#8�d��,`>mhY��; ���$�#����.��*���i��f�5������kT]k>JV�h��3���	 S��Y�{^�
��}��:tsm��ͤ8�0=f?C���n�L
0BǢ:Ty�b]:�X�0���CxZ��>{��%�vvܧ�s SŞs����)�!���y-�x�Uq���C�}O+s�':�t��w8J?��.�*.��Fu=tMM�r�yC�p�*С��"�(�B)O�{�b�߇o9�]�6z�]�� �N ������OA)��:9��e̺�"6a#@���^U��&ɛ7����=���,mk	HU	�u|�H-'��'uac?�D6(My�2�v�����<4.'8��, �Qm�u�h�� 8<u&�r1�_��������Y���U�農X͢�����=��A��z��6��<n����f 	p�� ��L��N��D	������i]48�C�]eh?�]_�uTi�X�����_�wE�j�}tm˜=���&�-�o7�`�AOE�T��k����h�	�~�}���`AO�h�꺁��S�f�֒ �����݄>tI%j���s�i[�Y�铷q	�%�U#��������.����ã��[W��l���@�
��t|B#�L���w���,���"\��]�?e�*'��޾�.����x>���p��]'6�3�#�z�
iA�;�Gχ;0�4��t@��|�]{zs1Vg)z���xق�X4G%�(��B\�#��q32g�C��Aͻy5���m#��BL��4t��?j*�%�	w`^d=F�XY�����m>�� �4ӊԸ�؆Ǐk{$����D�����Ro�NS��:RO]ݫt�����@5��h��)2��  ���jv3�������]�U#�k[�x� ��.za�E��ѣ�q�T3�A��^%�*(�;���vD�o��X�eI�ɪ� �tWQl����Zw�R�Py�%hQ�Ovs�ݠA>�K�P=�{�+{��Ɔ���۲���$ ��9���A�Ჷ�����	z�pdH�v�C����OǯD��=����Z��� >�\"\��0�X��"d2��*=�򫸂��ZM��2��^.�������TR� xI�ŗT����T���>���	��~����)�|��Ho9�4v�WW������T���(��z�\�����K��{�B �V�����.�j��B����JM	��<D9{���ă�b���Ϋ�?�s�7@��f;3&�OW�8�uJE	�Ԣ���ro�a��J��h��+�a-���o9e,\VOu�^�"�Ǿ��1��,�VW���ۃ���8�U����7��_�k�qޭq�ؘ�w�2�jzxh �v9�9��dǚ"[M�[�<0p�^��^w�������?��v�`�9R�?Z��Z��bC4��+���������S�F������K�9�cɀff^+"]��Ž5	���D3���c������¸L�u�/��E��!M�W���W	��_w�{�ǔ1$:�� ���k_x��v�4�8�v�ȅh9�n���������m]�z���Ɠ�ڋ��-ZI��L���T����L�1�1sk�W&�U������+��G+�q����1�B�N�ӵ�H�˜��Xt	�.@�]�4�2<J��Ƈ�l���U ��o�l{�?t��o�aW������?"��;Q1�Yx���� �$�FM�E�1:��
��S�� >�D��t�E{/~���.I'�C����j���'������\��]�"��!�A�V�M���[Um��5@$��u[a�1�j����e^-�,4!��1N#<���\C	���.���|]���fC�I^0���.��}���/g䪱%.U��Q�p��v���V.�:��:��J,ݣEn��6��}/5 uN�7rW�.�"��z��M�����ޅ|f�>XJ]��2�s���c�Cpo��2��6����>I���>�|�;�#zR���X�K����'$������1�B��$ŵ�&��3t��(�K�8S���q�������ޅ�ܕ��c�T��8B?̾Y��y�{���f|�,z}��8��M�"��Eq�>ݞ��z�~�gh�v���ͼ-tF�ZD�t�n
�g�$��U���c���Gy�l�zӢ�`��t�w7:�r{k ��8��W��>�s2����9h����%���M�ъ��F_��m$L��-�e˳�����z)��H��Q\A\��,�g?ǜ�7�i��s�(�etܒ�5�����)���l��F�DC5�{}��������1,�J��2���RG)j݌+x�F�0C�8;�)��+xn��p��(�Y��*��3x��,�]��A�'흝����O���(s��¿OV�W|�x�&��A.��ˡ��v?�1	7��s���'Q	wc=��LN��_���B�}�r�g�2Sz"a��͠��<�3Q�4[E�d3�hk��osO��Ϋ�A��ߓyQ1sx��~)z�������w�Y��ȧ���H���?tt�/@�(�@�oekH��N�`�4�4��
�Y
��;(g�O�Sy���j�����ST�!h���\	��H��gv�C���/��ǧL��#\A<	 ��Q9��%�d1�7 �%�wJyz��`�E|�o�� h����,��C�?1{Pb��
i�d��po�~���p; �s~��z�]\W� �]��owe�bmf��j��H��u�tu��X�ZҶ�Ƥ�Y0�Nj �]/T��}���`(G���C�_L�Ŀ�A���}B�T�]�Ʌ+Pl��lx��$��L�`�.fS1�^.��Ό�?�̍ρG\�^L��K==o4+(��W�`�]e�?��� � �'���\n=Xu��WO�M����(��`B��ms�!a�����a���GU�d]H�?�xk������7޹�o�6Mt���h��W��Z�e�/�7���v��&�n�&�£;4�sR�� �� �Z�Z4�:3�{��I������i�p"���c�# Z��W���9��P��D	�Z5�>)�1j�R�o��_�mi�>V�T�IJO�����o;���_�8��9�*�;�J���?��#�I�Yx�|ޠ��aqU�e�Qv���Zq �����0�Uz<�a2�j7��R��*~V�.��@�se�|J�5*����}*|��x�����'�R����ePs��̌���ypPo2����uj47+�#� �Ճ.'oG����~E���K����x{���(�L�9y��3 �ܾ��e���g��+>��l��m�[��U�����/bf��R���P�yI��1v�򵰏V�/1�v�slDB8�C��:�j�]*Ǜ�q�pK'z�҇�r�k��䵇�}ȟc)W��;��i缍[�l1�NG0��K��LF�[��pxi8���eEK;[���� �Jq{}�j�Ja����Ըt/&/�);��[	��-7��烓��@�G�G��j��`@�J�z'$M*d��YBW���߉���*���a�'�D��_�k���D'�h����ݨ;�����b�2�РNWp��,5�o�1՛}B({Ӿ��l����D��e�ш<|
�V�8@=yfk��$�'�S��
'�Y��WJ��s��P���jo���*��i��@r:�Ќ��O�<��t��� w��8vQ�X�4�� @�N���1�ZG�T���#��j���p-#O�[�q�I�3$�*�D�KuS��;qU�%��6�	 Vh�������U�.�R�`Kv��ҵ�#��^>#]:W�F�E�������b���0���x�Zw�oǋ�Wh�ӻhx����o F�s��H�����,��"�=ZwKR��C�\v%��� Y"8��-����M�E�ȾN6��E�T�2�I--�Dm�"s�*soЩYe������#�, �����Y������諫�ρ�-�Z�|�2�26*[X��5Y���@R�5�v֝��0���vj�h��eZAL��T�5�NRsZ����U�����1���%@��ꐹIe^Vr�+}W@�G�nV	.�NbwV]Ѭ�'e�=��  �$:���5~��7�LŬ��1"f ��y���h][;��w`G�>�� ��v�x�Y�d@�8r�H!��7��`}'��5s�g�;�q?��l�)��h���׊����7��W��ʷ�J��
�n%�1/�o��1q��[�����]W��v��M�{��O�ς`t�P�3����?�����tGP���'��rxz��o㥝���bx����x��|Q��M3y�� ��>��� o�?i?����C������ �^f�m��N�*�H6�_�0����,��2�H�-M��J�~A�\�M#�6z�!����,��?�ॹ�0�m0(@�Ö���{҆�E��2�k� a ׯE�0�����oA7����1��P)�&�&/vڰR���@�4L.���pW��+o��Q�	�=��Qu2�C�8������ȩ����l	�߇�u���O��+^�#.~b���	�80�����k����Q�w!���ʵ��PC�{(<r�e�5i����w��澋��f����#B�WA�����/��4�ek�&E�rzJv}�8n2��>��m���ڣ�.e�%^����BQ:�Ig5j�Hm�Y.קdz��ރ���%F��l�E|���3x/:?���?�A��L<�k1�)�_����C�!%�Ex;�L]��>{�z��V��k<L�~L��2$6JdӲ�	F�^�\|BrJ�p��M��[]`˴G�bA���U�"�M�Buq�N)�SO!� ���!�)�x�a5�x�̎_C�#�q���?�� �P{�YV�6o����!�s�t��RH��0\i8�;��u+ȕ�=(K�zyGM���9Rf�$=��I@�rm�ZԺTLJu�!~LWɶ�ӄ:F���!ɋ��C<����)P�������MȌ�	�U���A�@�N�����NlaBl�9�*7�k�Ϛ����.�k�^��׀��>D�x�I2_d7��lr�#�(M��m-���թ���ܓ}�z8�Q�@7bl4�5Fu�kQU�];ݟ=��0�H��b{��N"g���!{|���'*{Q�T�A<��J!Df Ou1�p�����;.��`m4߯�sy����{�B�PZ�Kl��d�]R�g�F\�T��y��I������@	�ѯ�����%���
g��;�g�:-G*�͸�t��&���� ����~l[~"���XN�pDHW6�M��x��?S(R�*��
��|��<��G��I���(��^��1��R���X�x@��W0�l~����+���w ��d?vɕ�j�R_8R���"���ú�������D,�0�$��	�,a�0D��T�nH�֖Ѹ�LQ��"�we�����)�Q	�lql�����BIr*zك��5�`3�( ���-"�z�/�1���L�7^d��O��&��B��j���p���FV��Ld� qP�k+��@Ԉ�Hę�������.�`�`&'�|�] HL/��h�cL
�ꈊ�+�AX��A=�'Z�`
N�9�����$��Iz0Vg(+V5�;ޏ]_�#��k���X�H X��8�ߑ�����Ü5n��i榞�ѐ��Iju��_��=X�EĀ�O��S+S�;��IȹX�H0�����~�J����.+��t�Px-���-�����n�z�ɔ��TJ�sl(�\�8�?/�\��ᶝ A!�Ny�� �q�Q�K�G�Y�XNOW_�kA9Y�^��^�g"��3��ް�uw�-K��w;���*m���C�ͩ���[oԄ�A�����|�Aj9)=yN&O�^��+��it:�8y��4�lM�|��uB��>���'/b�%@2���ς�~�����K��G�����/��v�R���~�e����3�^#.\Q�"=r�c>Y�2(������L�)�RZP��ӁY 5��]�QS�:�Ƞ�9��H��;�����K����P��iXF���ݍK��	�QY?���2���h�i��&.6�K<6?ę�R]9v� �!#X`e�鄘Y�-��"m����.�_��E��L]y T��Wn����M����J!B�� �}Ϛ}���e�ʒ*�ؗc0�dg$�m�[���{�,���ߙ�<���<�{�{R�Y�W�'�e`��_3ƨ2T�#��{Y�A�8G�8�(ѥW�}S>�<	?oJ���K��g������kod���}��'/g���O�.�"@������9V[�5`��M���2 �̄�e�\��Xߑn��r�O�n�o��R}�}4��n�g&+*j�3�\m\� .Ȋ�;x�P�'�M�������F=��*P���Y�)�L((�	�� ;!�l�b�+�W 4v9����1���;M��f:=74�XNw*�{X��?uC�U��$�GrobH]C1�Gw~Gf=��h�!�G�(>�n�>}�J#&4�2�o��v��,]�8d�S�?L�r\��gCլ�_�����S��:��h׋��	��e����v��S@V��C�}�������o-�U�W%�'T����v�юO�UĬ��_��E)��ۻG,^���g�w��6�y�	PL���6le_��R������"�w�)s�'i��kb��a��﬉��`���f�c��0������
�
qHD��Gt�M��.�k����3w�{�3�:��K1��.�2�ك�:B��z`�m�rS�(@:�0+����W�lI����n� ��>��u�S����5�t�k˟g��eÚo�]�,��ה7,�o�����zA:�(.<h�3��墣�E�_�>�������g��]�ډ[ty��_#S����my.�& i=` kh�\ս���BnۦO ]8	�IF<qg��还<-��VS8]c	����?�^����	0�� q2 $ׄ����Nx�ó~�Sp�O�9q�����h�_<gW�|�Bp{��%tbn�N�ȡ[�]�@Г����&'�u��D����������f�Dz;���O��<d6���~��1��T`��ob%���h�S�f�*��Y��̀@l��qn}	�?����?�t��'���1�n a�7����+o�N<�M��1苒!`���V-��o��՛o�T��캫8b!�n��6=���?V��0�*P	\c j��*���g�\5X�V|l0S��$��]:߹`E�������E}I�R�(4(������[��-c�y���"(�X҅�����E^î(�ѻK��+��_��������Lx��~�rk��N�0�䭁��;��6�_�/�< ^Ȗ��:|yK���Y��`Axp��&�?ua��4�pJQ�����	��@�p˺z-s�?-/���egt]�}�+��wf��Y�Mp!vg�/�jj�J6�15	1zg�����-�ٽ�<	b�?i�4�5^���U����`<�fy|��mP��U���6�0�	n׫Q�x��a�����1A����A
�H���B<Th'e�ډ;�t�?��GН/	ӿA;_sh����݇�;?}�[4��{'��k�1:z��
�"e�7�m���@D3�T���{�H�`
k
^՝� �'y�4<rwpu~Յ�`2{ uee���hg��|t�\�t����2�C�Ԑt�b
��^�D	�!y�.��p�{
��.g�R�cU�-������ۑ�y�#?�KM�Z2�駘��Z@J)V�\��=�{0(�ï�*�������Q���z�t���|�.?��ea]��p(�	�3[��:�Hh���	�[��(	�~�^�ⅴ��������Lg�H�6�a��kW��Ar5�-Y��L��y���FPp���f�nhɱ����T�Z��o��~^-!��Z�S��`UP�ϭ9�֡���K�&�������1���@xѮm1�n?�s����h;��� �J.�ܖ�O�l �z�5Y�8�u������0�?��Z�etN���i$�\�	�Nm����6�8x׉�BM�w�JѰ1`0�KW�:H4�Nlm7W~E{70�}O����0��	!in-�O��;�)	o��J�f�LR}z	/����4ޣ����(Eð6`'��E�0�S�㒥�]k��.��<�+_�$2�Mg����A��:K�+�x�@��G���q��-�'���%z:�t�(�>@ eiZ��nd���|j�8��z_g�/�i+Cr����4�(���<�&�3� �p!��kp>t]�P��#Q�
@Iç&�,k��p�T=�cP�=H*Y�$���P!�����U$s~�5e1e�Q&���Y���͙4����럿<��x���s5��O����G}9��{�����''�+����>����W��Y;'�&�8?��B��mɈ1��|7�P�p�_"C�6;���_{{��w����:N+Z���>L�?>�q�j�e=���a�z̴p�|�|�~��1>�g���>�xtr��	tu�S��?����:�P�k�|��l�c9�kS��I�;��dA-�n�>=i�=od��z�,�͖�1�j���\��8U�s��>��p��^�Ì!��:��|&t�LV�!\���ӴP�8��q�L��7,l4{���S��p9W4=k�WR7F����: t���Um�8y�뾧���0-߫u�9�jb�㏤®�M�A!)�"�i}���ۏ��x�&�i�38G�q㫨:�
�|�Ęf��q���О�*��AT��I�!��Όxbg٧~�l\ �|6{�@>!c{jpJ�U`=o7ae�'~��PPdx��@���� ��oo���L�
�D;����D5gٱ3��A�ί'�z�J} �FL{�9�)#cB�-i���E��AY��O��W�����������gB�s�mm88���a.�f̺��1<\_L����5���y�Q�������1�tl�9�q��� �%�:}f:��3(F�*.��i����;�Omr��M���LI-�� l�	���v_�C�N�u��B��0l�����O-��U��Ni�֛I�嚴#��c���>f�u��E^�>?��J��ar��o��"�QS'��Qm,�~��?c��D�~SU�C�eO��\1��Iiȟ��䞏�M=rVrȮ #q���������ͦ�M^���M�F���_gb��Ͼ��Tj�p��+��_�{@l���Gڥn��e;<�W͘O�����4��z"?�C��P�cU����ZgĜ/�����[�^�V�˶<[�X�<7T����Q���:�|��d��i	��Z�î�#��}f��=��9n��������{Fz�9Jg�����	�U�h���W��N��d�T_�x��jd&�̨-W����Ji�3i�%g��9�1�����6e<����t[I���,σ�n�釅@tY�co�˗���)�YL����yǢ�5i��Bx��@|+����'+ +#�̕�Yd7Z�*�Hg��L�د3+Ε��AH-�*��C9C_�t�cj�UB��'����1�=�% %�� �^��퐳\�_����M�}����T�]���+�"V��ES�$'���;*fB8���	�7|��:~M-V�������VN��O�!#+l��2�f�������:�a���,,r&{~a��b��gw��ȉ՞�z���z���@������%O�N� ��}�/�	D�! �M�d�/��~eǙ�Z�q�i�3�?�Ƕ�ݼ����V��U����@b��(�W�w/�/{�o"t���=�IQ���*8��+�
�-���#5$���oVlu3����U�����h��ح~�������gߊ�iٗq��ᩯ�5��jo|��4Y�}�e���L�t���M`�/�UѼ��N�<	f	��!�1 Fq�I���IK����:VXY��~u�v+?�&����V�.�נ��l
F=��i�5"M��/b� \)�+����S{�n�O���k�~�bZ&Y�����x]�o���۫?����Tbh��`�kZ*�@���4б���"��}�X��U��Y(���a�K�vU��8����X~��ɡ�:|�2�AV:�.�)�KJ�����+��QǘX��j��ט��B0�v�%ݔX����zI�����1�>I�*v��N:�T�S�>��}Fc��~�G�d��Q�U�,�m�O�,\ɯ}A>�My�r	4X��M�|��}�.~������䳎�UA\�/�>ԑ��w�v\��3$�֥%�3�Fa�%��tII�2��a�b��6���,�=?㱬r�-"22�#%�����m�.4�_�2���|e"����\_@/��������C�d��C���ȴ$�۵��{�8���Z��dx>����9����ۼ�;��2ۖb��HǬg����Mj��#���(lE�^pm_6��шL*�(40�W�ǯ�=�/�"K^����?Ȏ�Q}�i�rQ���r�Ja��pJ(E(�O�èˤ���?j��tɻ*1�3CQ�ǙV�f�Xe�7����4X�M��zm��N�;1A$��X��=�L����h$^'hB�j
 A���+%I�X��£}D/dl�,�j[tPRHB�N��u�9�l�����1����4�_����ev�o�D���P$�PXL���ZiJQL����Tr|�;���1Ӫ�e.�-�d��7�S�6�Tj�s#u`�a^Y	��o��va��<�5�~��Г�	�L�E�\�a�W�D���ݶ�M�g��P\c�,-�أX�ƚ)��`��!/\#���wC��Ċ ����eb=��<*�-cp
td�u?ɕvO�N���v�1�jgEmyE(���\��a��G�Ω_�Hˇ�v�
�X
n9�hj9�I��5Q�z�l��5���>�j��A}Q�0�j+�O��PjȆ����Ga�����#֑��s�5��$�7}C�"b&�Ol��'
�DՏC1�� �j��C�l�uGd��{����8x� ��z6	��nTc�ρ qr�k��ZJ�5X��A%�=)���}����ȩ� p�c�rn[�v�8n�j^�@���`^Y�3pxe}��ez�1����Bmi�֛q6���)�я�g���G�+j�}!���aixW 1�Vj��m��z��Ї���,)i�1��k�JdW�
;&��m�Ѯ�l_6KE���yX��x�v�����2�p�\�A潸��P�\˩��G}ɳ�Qli��m'��p�E��хGNj��f��e�j���1�fim�� �T8��O�E����˿�6П���B��q�='��������
!Q7E�4h�b��e�Qf�Sb��D	�� �J�m�hj�Ciq�����\�t�3���6��H�l�� V�c�m�DK���:�]�i>G�L��^��_Cy����v�L.�L~t�K��Ӈ�g�t�C2��!g��sdK�*j=3/�*1;L��<��=:�|��)m���4@�����"W\'h����-���{���c�y.�9��d��緋wTeM^H��Ik�m"{�����ph=Ym��ǩ~���yD���L#9Z[}�z�����y�W&CE��u�O����-�.�pð�/�N���HG��N�~�$r������%2 ��0o����C�B�|+ef���8��L�J ��7Yq���t��om^6�K}�>wO�X�jq�_(�z�X<�@"�C|5��d*�rl�E��[��ֵ����$���:C3��X�z�F��d�<Gy^'���L���
]]3Ɨ`1��GTo���2���w�e�hY�>/��^&����CGHA��1��&��9�.�e���B?mZ�cnS�����P��,ʮx�Gm�yMh���%��n�d�Q�,����/��h<q�ʹ�+nbO������1�L��e�-��|<4��a������@3�n5^w��o��PQ���f���ōt�?�s�:HKvf��y�2��M�1�$���ǝq2��qg����W��'lфTӇ���Ss�x��v9�cL>r��/S���W?��Ƕ��C�#�_=�G��;�=(&V�>={#�E¼�=Zb_�L}���UB��j��x��$����6A~�Q��K��ݩg[�dU�Si�9���w,4s�"�������D&�k�μ!�-�'����\ӾE%�.� FG*&�r?o6?��Jv��ު�3A����x��k��{4P?�ߝlm�T��.bF"��:F�L2�:�st�Q]���T)w���@S�T��u*H���//߁^�Ψ�@�b<�e1�>���F5�U��=C����p����+A5���bk���*��⯳�pn��H]۵���N"�;7��dq+Rܫ�6gM*���M�9�s�,�$�A�+�fW�_�-<�?���P��t�C�N�=�a��|�6i���׽�u�m�0>"["͔������Wvg�P=ƽC�L%�%7��G��Z�=��v��v�h�;;)�٤��0�T��C֬������᱁ý]ب�y���_�ɱ�ԯ͒�{�����[+=	���p�%�)����Q{��b{���F����c��&n6w��� AXZ9�]�ܝ^�p�}C}���.���}�$/BE��͊d�� �5ȟ7.ܩ��� Hʼ,��[��[C�-�(�P����QQ�)�G�#�UpqJų��s�����k9mI�^_�]�b�l�iz%h��]���)�BYH�[�X�ZɄ�o�Ou���/�"�"�����3��,��}'�����{`�u5��H}��"�ӽ���%��||��	.�C��	�3?��h`B>� "�5O�;4�����A�iiE��)D1|@�i�=�p�^_������̓[L-4��5�@��F�)���ZKm|3Pf�"�ƟR�q��8��!�V�*�� 9#���G}XQМ>��$j�^K��B�xh}b�g��B=���A�.�����Hi��������_�`���Fk�,��@�#w��c�m��ڴ�7}�2l�׽l�!eفY��$Z�>a��S�w B�nY!禱IY�qNw���c��HM�r��#S{�M��ų�Xj5�t�������Ƹ*��$"���B ��C�#-D��s��߉��h��0h� ��>�R�����>�Ǧ/ u�o+�%C��.�dD6�����ѕ��G��H�(�ٿ*��v�b����l�+R���W7�e�\���OC�>"���([j�|תM��+BN�յy�#�2�Nc���+S��q��0�3oS>�Wz�Ω��'�A�A�K�k��G�����6dۢ�_ H��n�W0�U��<�Ed���@�[��WJ![P����ق-=�����X���U�qd�X�Cg�؞a�}oӾ�;��ˀ7.��
v�t�v|_.�@�=b̆v_LJD:U�����mg��&�O�(��2S��UEEA��n�|���ǳ?I-ͯ/����ۘ}��ez״�ќ�����N4}�J&VH��f���jB���i%�a���4\5�����Y"[E*�V��v�Tr���36��/�����DB������P0�a?Ud	;U�%^��U���d���m�� ~��?i�&d��k��IHĩf���31t�P΀����[�Mb���ČeS�3�ڵ�~�}�4�xa��GbS���Դ��~��b\����QAվ;��Q�5Cu���9o��ۇ���C�~�5G'[����m�H�A���6�瘫!���ؿ�Z&ܸ��?-�B�ߧ���g��>9@���BJ}/3����D/�2�e����U3�f��Z��1^au�gO�i�B.:���[~
��;#�9i�Q!YN��ъ�U(�����K�r�/T�^���)��<���������V��[�����P�$^R�Z�{I@��p��jc1D�t�r�!i�8v�*�y������ït.u�;���!�� ��N�P�"vIqo=_f���qE�wZNI{�$�FP�C��[���y�l�K{=mտ�I���9J�"���G?z��}���Ї
v��2�F��\F�Л�9Ax�l �� ��Dñgg<�KwK���wv_@����n� �HL�c�]3���"���뭂�)}�bEHDo)��[�Ib$����X�uGsbg����<!rd����q�)u0��]w3�8��(�@����#�(w;��9v���Bz����X2;�8��7�6�� ��r n��T7-�˷�
��"U��Gdn,�x�ch"f��{3�>�Y��*}P�3�%���)Q'��JG�*ʢ`�/������M)�K; S,ӿ �a�[�����qo�>��x�A��K�gV��z��G
ެe9�_L>,���E�#����n��o���I�]h���ta}����Y�i�_5� %�ώI��Oj>�8G�=��6����_��C�By-D�6DoY�P��u�`��QԀ�'r��mE)��1����jn;����9|��@�b����3����M�,|�K1N�Gm~s�R�'2^�{�&�Ɋ>���&Z�0�k��t������C�g���G���QŗE�*v*!���ߟP8a�];H�<����섾^;�:$W+K�CzQ�!ȱGn�ʗ݄�vi�����}@�Ї)bh*1�h�����]#��p��1r`O"F�0K�b��ΠfHi2G|�Y�A�D��	Pg��p�����>�]-�Y�~��A����HI�t�9������}�Wq[gS	p�"/J,�k;�u/a��<.���������`1���� ՆNh����<�ne�\���D��C��
J����ں�N�/�v��AoL��LA�|]�R��ϋ�,�JK�j?�N���R�N�:���}W�h�- ye�������< ��m�$'+UYJj�e�=���ߨg��2�A7��R�����G��U ,b4:��A�+A�n� ]���W@S~Hi^�2�
�"��N�hS��2���"NAh4>�u�aS}˺�s:Z�XDN�7�$sq�w��
�Č0ƪ��;EB��"�oD[���leB�c̑�[�:�"�[��������ي8[F��ɐ�����٣mx�d���L����J�_�g�����1Ǆ������LG_-!:#}m"�+i�C��RMx�o5���=�'E�C(�.|�1�yDD6��Z0�����h!k��Mo�"��Q��Fj߷�������9�+�D��}�����e�^2dH�/�q�XW�U�횐�Q��:A�}���ŋBAp��$\���n�X����k�k�1y����"�s�"	�����	%���1�[y��@⛪�v�`�:�s*� �:J�\��s(�IF٪Э�1�#���Dg�1��x�KǄ�g��ԙ��	�I�b�	�-��2<�d�qu���J��ߧ;B�4\����،�!;���g7g�xa���%�_@[��w`^���
��Whji<�U�&#�m�5�&���Y���˼�tH�����!��w�(�뭢
.n����D(@�c�M~����z�c�>�$q��h�� ��	��a�gw�f/hy����$�B]��V����P$�����-_��)���b~��BYȬ�Q&��b�Ɲfs��R)�l�gg�^�����@����~S��=n�I�t[H���ǴP�R���-6K�#ᒋ-��S�i��v|4,~k;���M��6�Y����ce�rip�kT�����2�I���?�~���p2�}��^�Q���N�1-��s�Y늆��e@��{>��|���hN�"�E�bapH��NaL���:V�C�_x�U�^�$�'��!nw$�ЇQ7�J�a͞OJ��4���7���Dy�I�Slc�c�z�	��"�)�DԀl�]��'�����b?֤��O�*Iv�8	:}��\�&[&X�f<0�N���Y\��+��술VWip.�d�9�$��� 2��m9I_��ֲ8T"U��H�Yv��}���n��ͺ�č���$�������
��5b�_���aq)x�W�	���[�;�W[۶�a����(������t��-�
��:#��㡍�$���o�*�{��%�;'���i�V4��>&�h��������	-��e&�Xd�7?[R�V&1��!Z ��Ic5ez�f�u��	�R���j2�]lK#Я	=!\��Q���e~�����T�-\��!U�nף�}�y�qX)T�l��.X�V�4�@YI��4Ў�R+�nuqг�*�@��<V�1�a�KJP`Q�
�cyj>�k=�����~dC����.�A ٴ'���Ss5� �+C�˧r[����9�=�3힕�٘D ��κ�1���j6��ٚc�a�0��2(	1!K�g+ ��èYc�����q�"F6NBʎ�#�h�B�,!�[%/|+/)n[��ɿdAF����j���Xw��]�԰�Q��"|)*����L_��[t��p)�?o6kH��W	���1���ٖ���MS����|���B�QQ9�,R�|��j�g''����_C�m8��˿�Ėm�(튓��m����+�Ti��> ~7q�`0c��]1v��_fz�o���x��9CeT���W&�*���wc�ب�n�e�$f��2]�5���)]K�8�OX�7�r��xh@5q��&j1l����PR<�=O���_k q��B�����Ҋ/���J��q�=coC���kX�4h���0���U�CyK/�5I".vfr�p�X��V6��]��ʷt��|_h�/h[�%�	��آѢ�'�
�	����9���TP!}cU�r?g�B�RY �9�WR����!��i��������'�o��ٿ:��g�0,�,0����~���|N	�yC9{�*�ԝ��w��ƙ����l?yX\��y��H�vA�����`G��o$���a��)g�������^�pZX���+z�q�g�� ����۱ק+���u7����]ö�{�B�X>2bܑ�q>$?]e�<�<g������I�����ߊT��2�+�oj�(�}�����z\R����������K��q�=�A�I�~��*���s���ǪE��}2}����H��#��٧���/�W�r�)��6̵���}V�q�����% �����CJ{��RV��(X����b@#ʏ����F9�:�t����s��W�Ӏ����Y��HG��o��`E �Zz
��pɁqL؁H�ed���D>��򼅡�D�<Gkc��"��*~Η�k^�GI��J�VȂ��H���,����xO�}��������c m�%:6`7����Q6��BA����߃5v�C�~	8��7}i�F+��o�zI�vB�ڜo�XQ�=�;u:m���ӗ�'[�F	X�^�GL1�E���}�>>k~����M�W�2ϵ�tE���đ�Hz�i�:��ev@0HK��qiY��MP��Tx�c�I�ŀ���oǊ��n|_�ϩ�e"�".;�\(S-<m�!�$���h�DG�J�*����nY��K�N���3}͡0��=��D����)�Z��2�%eq�`��>�]0�Q��"���Sp�*��ZŘ��,F�'�ڙ�^i��b^����!,, X���] ��Y�S�;r��n���̵��B&��@jW�.���1�Y�i{��1ot#�~N�>gA��,Y|�k��ޣ�A�F�f�:i�Е���:�:�q߳ϣ�K�5�3�[:D��t��������������vC
擔L�%Z����-���N'�_�♟�Z\�S�� ?�P���	hb�i��������sdd������;���L�j(���gDT�d�%�q	-�����Ľ �1�vΥBS��T�/}{Hy]c�n��=��v#���%����6[>58#�  ڵ~B"�n��g��� �܄c�r,����
C/�pR:�L�V�j��p��V �=V�Ozɺ��C/?��Q��By�\��|ؑ��_R�rYk���b���GS�u����J�_�����_Ĥ�K=�����:ǃƶ��{[��-������Vgق���d��w �$m'�(�����P��d&�*�+ŵ.t���^I�ZUü��5�!�*�A>�U���>�ƅ��U�vLCh�G��)�הּ����9_�۝�8�_�@��u�ݚ���s�}�&�0�k�w��#E�4���_�� ����.w�K*���?��޽=S�aϽ�#�(�թe���Uآ������|~u��ؓ��F(��+0�����a�F�o��cJ^�ǳ�N te�;�g9(��� ��R�b�N.��u?�7�N���C��T���F�k|�r�X1���_�?��"�L�P��*/|,[d%������#p�s��k��D�s�rSÔ�(����7a�Q���לk��%$N,�Ś�r�Gw��!/�Y�i�>��Oճal-��h��\ާnG���#��qk���2s%��;kg��y~�R��&d�+��n�������;~D�6�\0���Gɧ`���ʴ,�����2�A�����9Z�,>��{��w� ���Uh�mK6�P�v�[�Bg�cS<���K{�j,�4/�}��0������cbJ�6q˓"����^/�i;�m�%B�[\� C�XD�a\�݉d�NUܱ2��4یM�ݵ�L���P0��jD�F���Bht���s�0'��v�bwp�qẵ��o�*��Fd���|c�H�u�uF�rvzW�5�YSp#�Z�qXM��?	0V�>Hx��;]Q���A�(��R�~�5^��I�6J"���Ä ���> u'x�Re�[I�C���Z��P��՘�*Ҕ��2�u-y�7ETR��D�����b!
�}�a:�9���@
�D���m���=yM�^�0>�lϽul���^�B�ږ��iC]��wE�Uz��Q��5�S�g�������n^���)��"b�N��cY͊�
0��k��/o�̉�9Y�L3��L�W�|}��I9�-Ő�������M>�n� �
L�y�O�d����e�Pt��S`����>��F�	��*'v`%�k���#<Y(e T��:!.]��{�v���굜��|�\{��	m.��$�1Y�e3r
򢏶�N�Z�t����0²���%G#f�v��_�*�$.ޞ�s����ZMŔ���f�l�?6�{?��p�U0����B3�#TUD��l�>����� ���s (�8.��%
YZ���4z̟�=��-it��`���ANA���J������Z�!�^G�|E>�J{�q%�F=�sX��a�3���ǯ DWT��}h2����8C�f�X�g���A`��=l��8�ȫH�����L������Z������@��ǆ)�,K�E�zU��
���r�f�WP���Mڅ�*�9����t5��#�t���X�� ;7�oӶ�j��B����#��7�ƃ�X݂���(B~CVR�����=����JnFO��?/y� �=�W����I��)hu�4�[�K�m��r�{Z�HM�$����$���e��.s�\˰��Z_@Y7@�����-�(�,�Ro���ۼ��T+��G�{d���]�xzv����8Q�A��}cX>�H��OO�Ee�6E"�67���	Nw�~�ٵYKG޶���iA�ǬU���e��\�b�?�X!5�VFl�S��_p;8�O=IK���l2\-#V��Tƥ�:�rtb�^q \�l��s�0C^�Z��J{� ?�"�$=���7��77Zo�U�I��+ϮC�M��a�k�6J�������-�,u>�"pE�	�H�۠¥h�,���v�qG��`�iU�~î�"��s�ۦ�8ϕB�5X�Z'����jϞ����J@S���"��S�������@ˌ������[ȋLg�:M��u��a��d�Kk���6`]��3����	X�Ut�_���]X�����7�4��#:��n98L(j�Ű���M��5�����Z�w�A��bh��5�!	o��yެ(m�� �1�S�8�$�1UB�(� G@�ܫ�ո0��;��,�h�dT+>J�L!���C6�ѭ>K�*r��`���b%�<I�\�/�����s�'NQ� �3z�38��=ӣ���oM�%?l��+��Kڏ=,ԗ�fls0l��g�lw��_ �v��
"�Zy��b���,��r�6q�p�n��� q#�Ǧ�xWeӱ,`����aRt���z�Ei�w�1!e(V P�t�Z;�ah��Ҽo5~FL��l�P
���Z��t�W6�$/㈶3��D���Y��`2��r��|���=J(�f��i�m�B���ew�+p-xN����4y\��+kV1��(��6l�*��+��Z��6;X�H��Kx�<G!n�B��2aW1]�v�1]q[�a�D5G��Ɉ�9��ĥ6�{��)�˺�� �����'<a������>f�i!D�L+��®��ԝt(/�Gsn� �'���7� B�3��e��2���uu�o��Ob�pki���CQ�Od�b�viN�ͺ�;�/+��;�_Z���u�H���܀��]���Q��#�f�j�[�3����8U˸�u�'S�
o�7�� xӻS�}��G��"q}�O���_<�,D��Łg�踞蘾���k�]E����*pbE>PZ &�bF�����<��FN�8M7�`u��hX�N�r���xpp�Yaǯ�=�Il{{o��cS�k�)öp��>��:�)�<�Vo4�s^A�!&n����{��AR.���b��94��/�
�w���յy@��B����^ML� ��kN3N?���0I<�L䖡��pc�+ ��k�W\m��еelE��Z^IP�XWoPRr�������#ׅ?�f���v�'����B�q�Y����7��W'���@;�w��.'G�s�j�E��4T���mi���[�d�1e[���~�j(K`W'�����?�j�@��!T��]d���gk�E��I]F���MJ:��o�`Ϧ+M�WQDg�7H��� +{v�i�8��]z��QE�b��ם�E�~x�[ �q��<�=���L�fY�7���}�t 
A�:A�-h����RM�B8�����}̔�%R���<��"Vܯ$x�1t�@ē^d`6��L�7|~W�V^���Ěݎ?Nu�� W�b�����"��
�g/����W����_?��Z���<��+���xqR-��v�����*aZ<N ��|VM+�w�� �Z;�Xc�%>����d�yu�k�|��/������3ٛ����=�g�GD����KB'l��y������d��^p!v��9��c���y��Y�
�&�=�RaGr�"$=׃S:ғ����>
L_�)�U1�W�m�<n����1'��%����$�������c�M�J�G�L�IOF]S�s�Վ�ή�C_����Z��NH�	� ,Y}�~.�w>
�haς-U�_ۣ�E׼a��3��P��D]dz������	<��W-�}O���ٺ�ū�����v;���.��M�j�G��z��p���vKH�����̈́6!H��rt��g����>e��!�{n=�jj	����Y�z�ќ_�Ni���l��I�w>6���f�޶�a	Y��{@��ݖ���oK���w������h�<~-ZZ'~��Ǐ#�1�r\˥7E%�]�r0�۹M���Y����r� N�z_Z���՘�*�+��!��M�u�.�fԿ��G�U\d�p�P�r'��������O���9�Z{�p8�u7��x���0���5�ϰ�B�ݿ���wuH)�6�a������٢G�mԨ.�kB���J,e`	�5�,�;z#0^�G%�YX��)��]�����vAX�Y��e�0��F�V22c�Pq�:Kg��+2�����#���G�O��'���?F�8�G*)Pn����%�qv>�-�lz�ױ�u��9v�h���tٍ��C߉�r�[�������v�\��35HB;
����>�ȹ {�kŁ�7d�>d��T	��T��$]ϓ۩�;/��p��WæWS�zm�"�$S>Q%B���_Ѵ�9��C"%Z� w`�ԡ�o�ߗ�&E�岅��	��2��JZ���*_�����;^���"�.�Vr�ʛ��"���>�	��8������P�@o���O�#:��!�7,t�ΣL�Đ*(�Q&*�����j�1?�/����t��<�`����`�!9]���E���y�G��oDy��xJ>�v{%�c���`3RZ�����c#{Q+��]�~��%ܒ�v��ݏ��n�T�B�^���p3�
K��2�v��V��d�)&���ծpA==�G?�
�sC��i��T��F>Z��NΆاr�=W[3���m��:a9vň�E�i�0�Mc��u[����ʽP�*�XM:�Pk�-���_�8E"w\��B�F*�n���b�!w�l�=�����w*b�ekD�B��|[��ey�E|M)8��7�G*�BDʨ��ĭ<���?�
F���p�*��k+�)St�U��t:|(�6��m)�O��E��Q+��o�H���\�����a]vkv.���W��n�危S��>�B�����F�%5�*��j�v�˳G�(��$E��P��0+{�Z��H�~5dϖ,��V@Tv?�v9}��UK�~�X�F�H�0��V���2Yb��*�#��@�:�_�Rx��^��7t������j��0|[��:���BC�evxʦ�D�r��� 6���kR��k"�ބ�M�������E�ŧk2��8Ŭ���6���\N.e6�D���[������u�\|E+�>��*o�V�k#s�8��WQ;�i�}h���j��\����s�UX*MT�ԿVm�rσ��1h���|�R�lz�G�F0��R]��ȴ��U#� sM�l����ل�2�~Z1�w0��T_��2g���8���(Ε;* *��_�.�jhR���D	��Ƌ��SX4����!�݈�=�c��#���y��S��k�}[�`O�>����!�=��W`N?��h��H/��V�Q�����Z"�ҥA �%/�|����A�x=�Y���^Z�zB��ZQE���d�#n��L~S����*T1t�ȼ��^��,��r,>?3q�ݧ4@����1���C�Ae��q�^����z>���~֛@�A�t��?�
DM�_ԙ�G�\�P��u�dg��m���óS��"��+d@��j?5�������˝������I��=�5a��2n��E��L�I��]u�W1�&m�ބQ���ա��R�Ϩ0���{�Ǭ$>(!��Я�Ɂt�O�<���.ZN�ui�5�::4LƆ���M/6i�`��s�u>��,ۯ����M:�N��W�`v!�К�8���Kat�ϣ� ,Z�~Ls�P��Dj��T�$��U��*}�As.���dI��hP�0�nx̝�V��$�bi��i�'�,�H@\�2��BhC��9�QjW[nqA�g������Ꝇ����m���Ra���y�":Ʉ�����3�a�y�ʽ�X/Q�n��b�sxD�P#�H4p�_���?��Ը�W���9����˭�)�T{�Q��N�4.x|�� �����Z�m14�炦�3 �J]�����(CŰ�=��]�V��;
�'΍���L��aE��(�ě��5?������j]fTk]�׸�M���N�����霿�X~�H�]�b��P�Y���$SP|�r4�2�[V�Q��[��܃|�7���P-������3��V�%�I�[0r�"-py�0�Gh�?Sm�(Ug ��1����þ���P�8S|I"��N��tS��:�j��{ R�~+K��]�n�ވ������7��Y���8O��"ﱘ��#u�<��Dܳ[�.���mmQ�;���\r�@B!��8�rV��[�|��|"�����5e؂s�S�m��	��܅j'�u��� 0�mo2.�l?���Q0��ћ/��rў��|�f�ݘgg)����~r�'h���kv�/��>����Rn^w'lL�:�G�ێ�g
��0)p�ͣǒ��ۼ:a!ʵw��M�<���$`��̻���ǜ�DfQ��Z@b4���焪�]y/���6�~᷅��0����Y����.�������aM�q�0���� AB���Fi%�%���"�5L@EEZ@@@B�ѣk�tw�Rb�6z4�k����7�q�Rw���'��y�, �A�'�d� 0��Euef3�ۏT��5x+�2_S�7�X�}77Wv�+���ϣ��8� ;TZ�r[�!�D�ʠ= �Q�����߂p'�޲BZ.�bCG�30ۖӖ9�ؚEb�j��F��	Z'ʅEG�8V{r7�O�W��We�Ǎ�O屚����p'Un�7Xi�u���Q(���
�n��&�}����b���h�?Ka�N��a��ɲ�5U~'Z��׻����M%��`L����見�pt#����ʏ����;�:�׈�Z��'��fO���1֨d������,�/��E��䷟cq���9�8�N���,��,�����7l���:�.P�f�S��ɗ��Hl=����G\	�x��a[�����?*#E]G��.�l���4�� �C��W����Z��y��G��.��.I�olZ�H����p�N#�c4QX���7(������P��667Q);4�I2�h���f(Z��5N����OI�f[y�����/m/]Z�"d7��4��$�7�E�<W�!o����G&�Y��]Eڣ�H���7�����2��+�V|�|N{(c]I'[GL��)���4l7��F}Ĳ|s���ϟɸ���7|�o��m�njT�ʋ��<$�xs�� K�2�{YIe�Η��r\PJ��G�t0�0i���\��%kv�9����b%��c b9�،ryA'{����͚-��[�N����R��]'�@f�vK��b��Ǥ�2о����ą	^�e	+����nE�v��$�6���V�����E����ƼT�У.��4�u���:[1�������C�㐛[^|�!H�)'G�E$�D.�����Yo������'�hRq(�.����鱣�q���\[6 H5/��Z{���6���@���PP�ˮ�~��Nt^̈���/���=�n��Y��L����ו�*yͥ�;�p�y��6��}��45�²�O�����]w�}����x6�Fk�����0+�L��i���h�}L?��4�i���V]ǀ|I���� Y����&&���noQ�)��x.]��ktj\K�:�g3�%�v( �~[��#y��	!�z/i�u-(7;��d8��8������;�׮_�c@9t��k��au~  ��_�~�&�/���F+�C�c _3��JqG��x���߻ͼ2���H/|y�	qy��zM�ʬ�	Er
k�e��N�'�iZu��S҄R�ٵI;\m����\�-����}(@%dc�R%��u�B����2Gj���/��O��R�2=����7�Q<�l��d>��n��I��[�� O�u�P]_bh34�N�s�'����w�Ls��a�Z�M.+�*�qV
1a��:�܉4��
@��jpWN����e������{Y.�I������ķ��@ꉓ���\j�N�ЩsKg�$[b�L*��P�����Q*�
ͩ�+�G�,�V�[WkU�F����z �Y�I��1E_$���X�9^�S��gRW� �%�H%dw�NG�,���O
��/g�2���y���h�P8�(��7�me���<����P�/ܽ�_�o54ЧW3n��������)R�߈!�CFA���X7N�5~
>2���/]A�N�Gw�m\����}ƙ�Hż���M9�mE��<Ù���%�n���]�z
�y�?d��u)N����p&�H/������a���;�o@��m�^0=���\`G
 �|hN�o� \3YQ,6��8�s�c$脸���@ƥ01I��^�0hԜ�X( í{�y�t�g��d_q��e����M�:�- �K�`�s��-N �d���Yp���]�����j��%>z�۔�@�_�&y��}��o��k֌���(���L&Q:���b��0�A���r���
��o�o��`s+�B�2�ʬH4���}�Υ����z!�e�����[�[��"���1����o蚵[I�N�R۝�n��e�R�Ӷ�X�tY1�ת�nf.҅%��v?����$^��L �� &@�̐�����*o��<�cJ�$�C��<�sA��`ho��)�ad��(B����-Z�13�> dv�_<Ox�OpA�
��3��]�a-�&��1%nya���\v���m��r�kYe�M��0�y\�ύ��=> ^��	hMO���z|��&�oIsV���>� 4$�FJR4��x̴8an�×�s6��AfO��Aqg������9:��z�T�$P�u��t9Ώ��i���Օ������a<]��ZW���K�L_s>����n,i��M��ҁ�[g_EB�_~&0�ˬqZצּjM�W����Fꦻo��~�:��ښ̳GF�C-{��A��?����X��xI
����2�K��ޱ/#�8+��B3�NB�4d�{��HU�C����z��	!��v�E@�(_{7q}��}nӷV��^��7�|�Lז-��4AML��3b��f�1V���s��Լ��d���,+�S1�I�p^_����+�c6X����GI���W ��c�71Z��q�|�0h�G�lÛBY����4^.e]����z��,�='��5Kb֢E���+~�Q�b�)�|Ҕ! 
�*6#��<=��X��i��9H��d��T�Q�����9����*��N�e��U`~��L�+������*t�x5l����]R�l��@Z�+�M����#%GW x��Բ������� ֽ$��"]���]0nkd����qYDcn�Ƃ��q��\ ����)�YUs���	��ly��^w�3Δ4�j�T�&�s'�L�f<5����,Ǿl���i�Ahn�[�ڭ)����.L�H[��5�/tfveo��Z��rqq�C���/2����3�:lv��!ɘ?��:C�
�t��d#76��'TCUR�N��Q��ܺ���餙R�6�֔17��ַ���P�%�M���inO���{�ي���'���	��3#����1V������0����2	��������O��˼(|�犙]F�m�ǖ�+���9�B��/�e��Y�.夏Q�vɯ����<�VwҒs�!�z� �]�ԯo�x�h-�[^a-q�4˚�on�ѧ����P�t�5��Z��&��g�Vb�G�FO̙��nY�v�Z�.�_�������q[]�%ճ���O-:� 43M�b�'����/4�%	��cc:��WF�i*H�п
�Rn�����?UX�I��S$%&��ݚ������<��;Ah�"� ْ��9�ka��ܠvw�)3{p�~�B�1�t���lI(`<���_m�Xr&2$:��-�A�zG�k֓0�<�Қ7G8N�%��lW`�ޙX(��H@�6�kP�j8��wRdtZ�ʺ�i��������%!R��idM��g�r{fۊ%1P�[�����V��c�VZݭ�e�����r0Г��y�hٽ����?t9<>��������GV��A8&0�[����`�j����볇<"�p{I�J ���g3�u&��������G�L��	��JV瀄�$zT�5��ޤ�E;�����K@�ON��`���AzP��q�c���}�W|���_|Z�1 �]���S�LFV�vT.J��o+����V�c�������-J}� ��2���-$?&�I� ܬ\���>�B�}�I�N���۽po�y�h��-��V��Qn��꜅R�#�+�ݠ���En��#b��K�����Zw�f��}cWrK�/D7k�(���[ķ���c���#��$��8:�N�X�LB��b�D`r�=�_�4=���̍�����w�\��].�100�E�i��J󅹢^Ӣ�c����=�,��m%��Vp(��xR��֒���OzY̋b�O�K+��|����t'4���*n� ��=n!���0�����(.Sq�S/���ˇ|�PXZ�d�k&��[�oہ-�5�~%��sY��� ��đ1�Wn9�F/t�j��F�����R�i���s-���0,��2�V��6�-Fiq��_����m5sE\g�D�eךq[�r��`MG��X�}#P����*��ԅ�Sr���*W�i��Cӳ� z�_`�}�PC�I�h��`.tz+�|��|��3?�F\/�(���}��������
jfQ	(%e�*�m��?(��@�$��Om�g�7j��u
��Gz.=�ta|2.P��v�Ί��::����"� �01�]g���R<����f�i�}+� ��W�	?3ӜXny�	�n�v�<��R$�"[<���x�W߲)�7����ʼN��7'L��H�]OY��;�Q�$hm�~�o��R�n/ǩb���]KD����%�~���ߐ��^��~��j%��Y���ڙ�ė^�Jѩ��A��Z�L#�$��w�C�;�$��8���x�h�-C�	Cͻ�����4> ����ٿ�����Y��म��e�󻓔I��i�8z�~��f_tLzϗb a�v��+���]��1+�s��6V���V@Q�-��<�ԣl]�|P��������B&[��%M+X:;;��O�<��E�z�,Eʿ�O<,��w�\(Π�[=�� �[�m�?����Y���k����n�G�}( aK�?���,2�Md�/
�o��&6,��X����(l�L�SYэ��h#�S��&}%B.漐�ч� ��O�[��ԯ2Q���OS��,���J�A�&�'+p�BbR(�>� ����|��$�\�m��x
�Q�,;ܷ�������j��c0d�l &�eg����l�s�^�l�d!��(�����5��U;2�H�FT��F�!O���-�WʝA#G�d��H�����B�WY����4�.��`=�d�="�y�*����$~<�Vd:ώLV�!��xb,��Mn������1'L��Q=L�9�דϱڑ�n*ja�a&=�_+4�.P$L��1%�	���5 
+��Y�l?2&�J]����ղ�;H��2wR�l�����X���� �������U� ��]�K�b��j�R� �O�fP�BHsJ��
˫p}*��C?d%���ߚ41��v
��w��	��B0� ����[5�V�)T-��
�w��K�eOG��$7�JT�ʚ�
J�YQ��ٹ�>���ϧ��]��q���}]�0�S�&ѽW���Ʀ�ye��DJ*7�a��߹݉�	��G����(�0�դ˖+/�@s*:���o)�X�'���bo�=�e]z֜�h�]����ų�R�Ν [y�F�pO�í;������;*6&r)X]6\�~��"&��ɭ[�f���ZsK1@��\$�٣%��t.��S��-�P5��*D������|�q5��z���<Lq���ۿ1Z2����?{��??��?��?m�3���?��&�O���w09go���vU����Z�4@1��^8���C�kd�M�hosJzdԴ�h��פ�v��"���8u#~I�'���7ˣ���Q�وl8w\�Q�	Wb�kk�q*�*�IqR�Å�O�8�i��w
��"�z ���t�E���zᵄ�BiW�|T�l\*S�����^|zv`�)�I:D��lF�Ccc��FY�D	���N���7~�a�¼��P�|
#`H��y/I���g�&��/�1O؇%��{��&󌢓dqO��wjaX�2.+���q�u c>��}��MGHOO���B^���	�F]�6��?P~���ˏ�}������������ū�/���*̈j��N�;��S5��Wi�U�h�I����%��)o$�X�'����x�^�Nj����6�Nw�;���wڼ�o�!�e�R	R�/�	zY�P��3<�Mi��5?v����J@o�\����&���n���K]��yi�w�s��Gȩ�����xj�n:	����Q�������!�ĽB���e�WuL��C����ֈ�M���Z�ư�H4�@�b�hg���g8ū��~7�V��^-#������Y#��J����q�$�:5�'z��nyL�yV�s���.�����<!�MW�I�q�g}%^�l_�65?!m)&t��=�5�^�ЉH���|9z8}��!Y��i||����㥕�+>����
�|��Ǭ��Fg���$ŉ��M��d�Kj��(���d�	�_��߇�+��xi]�5��������'h����mi/����;+E:����;d6}�s�XB���X���ǅm'�2�ʘ��5"��>�2��5�]S]k��V
�ʖ����G��<n�?{�z}6H��m����^!�v:�r^z��6kz��o{f����������Z��uf}�{�n�eXn&wSg�ɬ�-�����ߛ�U�m�Bb� �q��VW���0���)���_B����Q�l��_W6��B���^�\�@ؘ)�-���TM����]5a��g���¢�?�������4F�g4����;�3�s�2�F��0�M29���p��g���d#	L0
�ZJ�z�v�(�m-�](I�(]d��I?�y�ڨ�s+������r}J/��`
_�Fڳ���Ò�C��9'OFݪ:_O.�u�w����k��Ĉ�wk�B�n��j]�`܍�移����(������JF�\i���1Lպ/j'�G�H� �R�jXu�G�pPP��x�&U3Y�/��~�Y3	�Ǩ�.��5@���}n�RQR=�X5"���M���afzz�*G�^<�me��w�dWݎސ�C|�;�����F'Ů{�0��w�O����?l+��ZcËC�mO��Ƕi>���A�mY!��^c%Y���C����;�S��پen�\	��H�閑�;Y_J2�X���E��TG��#\������V[D���a-�&�m5g���u�O����
ɓ�x�y��N��Y�Ě%��n�|��ɕ(��� ?���*&Щ�>c��N}���~%>~�A�vy�i�	�L5�������'����YbM���\��XEe0�@�銕�I�Y���"�$<ݵ"F0 ��_����R�
�tEFDn>��f�M�L=M=�_�'į�@u���"���vv;+�&�`��Q���/�h�>!�7���Ք��ƣ*�����s�Qq<��%�U���1];2?����s=3ٻr�qn�(;���n��DH���m��"�:L=�0������w61"�-�����Jt����������8��d;<����~��i�Kn9Ϟ�[[~�ͻ��@Y�:it���D����'�:N6kw���
� P-
����w���io<�� DD��s�J�n���,��R�A?">n�����w.��9��?�S�/H��Y;Eo��ڌ���H �	���'��%��*++M���`=��`o���u��TF㶐0���Vꑗ���9)U�C�^ 㝰�ۢ35�W����9Hk�d�AO�B/��s�n=m�/j��mc��/�M�2u�\]���N��R=�Y�h?}��&v<�����x�N�.���hJ5f�/o�Z=� ���BM����z!J51i;!ȎeQ+���zi�CާGĒ�(F2���4D`�t˱!���З���|�3SU4B�t���w��K� d�nVڣ/�.{i��5	��K:���H�u4�x�n􎽛����O<��Y����=|�Ϧ|+���
��O��b�gC���-�9@��U7I�R�Y(� �^����!��䯺P�e�y\S�%�x�G<��8�zlydtnEd�&�4��T53 k�e5'>䓥�>�c����ǈ��e��V������m������^P�M���_f�a��1�ⰶ_�Ny]��L6r���ن<G;?|ć� n�`nЍ�~�頋�I.�+C���l��R�pPf�������g��<5'I2'
�c�)an�Ӝ����pW�b��~YV�<��2O��z&?��S�єQC-�CL�N�W[LXf`
����߈��>��&�N�ƒ�"�*�HD��%4���'-��o"��yOޢ���@��2qj����Ù�Bi�h�Zb6Y�sB�	@�����U���,���dW�R6Ά��P��7T��;�,=�I'�ꏭgl'3��ݺ�����WHYs��[��a��@��Eܼ4��{c�	�+�M��cN'��y�&u�%-�����Y�{ߊ�Y�{k����8^�o�=�A6�CT�d���P�7:s���
!��	���1ʐxu���X���9��wyו��*�6~������꟝�.s��G�\1:0� ��E�	��Ց$�	�0�2�����ɔX���6x�q����	UF��%�8������W�Wq.-W�Y����>�g�P���] w��>,��.�v�RU9�_��{��� �x`P���Bwc���P!_^R���]��k!�nrSD��*�=���.O>��߉�Ъ�6�L���۴BJ�-�%�m� �Z�T�5R���P��݈NU
P�T䇄>�	ںR@H"zq�^�č� \�>����^e�1+c��XK��#}� iXR��G3�V
MO�f��z�T'u��Ub�U��ah����bdp�D�b��@��'��R����C�O�5s���۾��|�c��}��j��6(�q)BT��+�+ �:�^V}S���7��$�G��ɞ�7�n��W�z�7j_��@(�6K{w�|�M��B�u��Tc+�d��v����r�<U�$�Di�׾��
����[��z�\��7i#3k�2|u�7� �@:��[wI�D�N�Ƿ(��ijNq�v�s�vh������W-����}�+׋ee�T���8�=y:�wFgFw�yK#�-�F����ǋO|�~��V�[,Õ!\�U�;/֙�@eWg� �}u���|���T0A]�����I�3��SE�n����b ���@�N/��Rq���A����^��j��8��H�1j���ݕd�fę�!^�H�%������a!,�#4ޏ`=��v���IW���[��|��4M�%�+S�թ	���7���>�H��z�'�7T�z�����-�(}F�N=��1��r�����-O��t<���v��p�LH0&�'��rמ����Z3�)�Qٻ���x��ʟ��q�d�K�>�i�5kO<�ȯ6u���{|�a��R�Nl��n�S+��@�N���� ��� ���Pҝ���ϐsX^yJEJw���.<�V3�:<a-C���U�Yȹ�S��י��vׯF�����<�N���W|�+��^P�J�����8{���r������ZAI-3��#<C��`r�tsep��O�p����)�BvFi�# q�H���i��h8YŠ��@?,ئ����_h4���u18h���d��r�)(e��8lU�9Z�H�}�WOl@=��|��������z!"ǳ�2t���P�T�k�v�B~��Y�ϗ����������(z��g�<�K�Od3��%�E��d��*_˜(���J��&Օ�OL����+���}�Le&��^��M��a� u Y7�����ȉ%U��W� R$�����-8�0���~d1ډ�X���.O�SQM{���}�CeH�ih�\���+����L;���g/�į�D��ao_�f�aK���������;m	<W"L���Vl��eK���[%iA�^��c#�4��B5f�L�r�� ���Xa�
���>��z��6_�r��hT%?�w.(��+�����[,�b~�Qf/�S��2{�l���XP������s�lQ9��ʿ���b���Uk�<>A͐hߕAٺ�3���X�V15OK��v�e�|7l��!���]Q��e��q�#��h/I�(
�ʳ��v8h7�&뾵��M��m��ҩ[O��%>�}c6)\���ڇ�o(�� J��ԇ�[��i��;P0���������fa�t����������z>�H*xĳ�
v�}����t�U1�ʛ(r���ؙg��2��<�4���w��C ��4������ظ?h�v��{6����q�t� �v�>��=o������pB��V�L�(Q��0���-m
�!T����<��K�M�3�s*_����ٽYI��+�h�-��>e"���!�
H�+$>$�G�*��$�2�3mJD�	P*z�D+��~wSs(2Ll\�Ob��o%����T��^�[N����):�#t&rC�k�y8��l�!i�,X���jl�p�:���/⥬W�֕&�]92�WH���С�������ʯ��1��fz��Gt�a���d���td<w'SN�-e��쫓��+c���0�?�́�?u�B���6Iv~�)<�b(.\���7}G��J$x�Q�4���͌+�v|��A����l���<1͸}�T�2��F�ke
 � �"���6��W�r�V�����~,�vZA���T���㇃?��գ%y��+V^>�-����H���Iq��a6���i׈8���rDs.Q f"Av�~�9�b��Y��R���� �D�d�i����^6�ꇜ_�Ĵ(��V�V]!���ʀ\�M�n
�<,��w#aBs��"�Sd�V���۫��<��!j��D���Uuԭ�k�:ϖ�F����]�Qv�/ʎ��Y��е_����'�d���p�ԕ���� -���}��RR1�r��z	���WH�!nᬺV��E$��sd��t2�����	$ͧ�'�����O���y��N���q�YߍY�&r���*�	��;�Hx�����XH�1�h��=��74��D=\����ưNȄ0K�Uu�$%�g��_)�T�fci8�E*�m��:��c,�^�PhLa���l��W9?�?�����2�8.?������ WNX�:E�W#2�Iyf��-`���8�Q���(��"'d;�.��ʍ�	�R'�P-Dq��7���6�ֲg|�t�����:.k�������z����"ɉ��S�u�5���^Z�Ffĩ���^�./��ҷ��M��H.�h|��0v/����F�j�.�����E���G�#����M"��J���B���qj��r�[�谄������'�5F�]�����>d���wo��6��u��z�M�@K��9�s�f����\D̘hqg*x�ü��Nd��P�n&��`�<�
��+Xq:�zY��U�؄GX�ˡߑ�+߈h���,J���f�1'F�Gx�H�Y��r���3������_�qs�t��o���RǠ�����G����Xm7�)���ߡA9M�h	,c���	4~�8���2��y��� `PV#���ZE �E����_�M#Mhq�1݈�����i~��$�,�!�j�����9_� ������y_�h�FG]�~Y�3�0J�=�7�q �'Y���W$������8�q%�0=�fPV�P����&��>��̚�iɛ|�W 'f�%/��V��0�g� �C��u1]P��ЗC���&�|ǹd�	w��Ɍ��xc'ٷ�>�0|z0*;sXu�������GXPX�8�e�i�]>9Rm�>(3!���{(UB�VJVMh��|��Ç
���7�����ml'��F���Ѷ�7�mT�"ؙ��p��O=�"�-�H���&��ec#��������?خ6�^F��6�9��4b&-	��>�$M�<����=rCf�P�FW�������p�c�����K�|	�}C?�"����y��PR�u"����?C�?C0
҉�d����un����{�-	�x�����o������%���9�q�p�9�i��'k��҂�s ]��H��% �چ�嗨��i*:�[��O��z��H}��a&�L%]iIW�*i`���]��Po��W)r�R�����d�a�}iO1��])E�����ϴf:�H�ry�iY�PԼ�gm���T�H-�z}�)�LW�Bv���4E��	@��"�*��_�.�����Y�aL���#��.f��9 �􎶰�T5q���! ���̵�U��Ab��: a�N={8G�Ӳ���*����e#��E���{}P~2x�}d/�4�-�,g;ԨR��]z��H�^�O�[C9s��N�}u��J�}Cƨ��UqiO%j� :f���0ᨤ�I�f��.)��%	e+m�i�Co�R~�涍s�8�S���dj�v�����Θ����W�N������D&�2v�Y�8�;�2{&63
�I�D���2��儐�,>�_G��9�z�k_F>�Q�.jk6T�,?��>c(���L�8
�E�b��ρe��/��;L�6w�15� �l����d��h��Glh/%:���;�k]Pk�eq�\|�'f�֦��iS0�����Ę�F� F�BT{����C����k�����і:��o�~.��\����0(���)<<:�UBڼ���C8�#v|u��h&6ˁ)�S�śo2���6����� Z}�r��mc��__	���G�_dN���cX�+'kj�B�ڹ�qҐ��C�p*�W���wM�*z?gWV� c�mm�Z�5:
8�`9�(�:B^Nc��]�C�Z��/e,S{�S�$f��oq��t'��Y@OǨgY֦�;�N﷟1�-3�+`<?5ew5���f{Y`�u]?}�*D٤7j2{����4�p_ٟ�^�T3������
�����b6뙏Y��LJ��E����?�*�ݰI�.��>|gӹ���3,b���A��"�W��?�l��nuў?�9�i���?i=��8kM黤`%�4�
� ѐ��#
���v���O㏗���L�,��lM�A�����>sIU��@!�*N)�j�6�(��Pl�I��į�u������̚:���A���K|��nj4����׾�����~��?��r�,8����Ė�%ę�R�v�����#�k�]�Z	����ᙡ5ΓP����D�ӧK��ok,|���#@oӎ 'X�Ϛ���t;�T�̗���l��$�#�+=�0�f6H��U�R�e# �������tm���q��X��v8c.�0�Q����Y�)&�*��i�XFY17ђW(�Z��{���Ͽ"f[{Qa����^4����V?�D�Tu���l�S�U��A���=#D~J�,��ĝ*���uL�'v�5{�1v8�'E �й2�<�)"b�m��ܲ;A�M6��Ӄ���u�d��b8��$A���P�u�$Rg�/z��Qy��sx���� t3�X4W��@ar.@넕-�G��o����N�+$��W��Ye;\O��`ɨ8���{�6V
�{���8��V�� E��8��4p��䥯*���CV�x���ȏ@�}pn�|�9��u?I�&]�BElCc΋Qb�Ү�u�{ŭDa�7�`@��������λ
 )���,��_
*7�����5�b-���ں�qGEO"#��h ���Zό��{��딕��.��5���kVg4x_!��$E�v.]v��
�+y��
����g����k$�e���Ws5���k���K��4x�P�ə�<�H��Gbq*zZ�9<ľՋqTW�ШBN}12Z�G|��k {�wՇK� �KC�m(V�/�7�n��ns�q.���d���x�=-��hd]�����d��h�B�zl����ߴ����8�Ei������ͭ,GR�)e�xU�N�mnOx�FoۮM�02�ڋWr�'�4��Īg��ǟ%rnZ��`�I�C��E7�9a͇���2����b/��ل+�~�Ò���"�}1���HB��U'�تP*56���d(��r��&�q'8/#u�\���g�$�D=�AD4�&57�3���s���w5o}S�90����P��*%�m�k||��&��L��|G����x묦���}��tz-ũ��oT�@�1�<0=�2u�S>�,�	4-���辚��%��,G�Q�(���t}�*&��P뗑�I���ȅ���u$���p< g��[&8�,� �O��7#�{u��)yr���\��C0>����{om����*��
���+�%߉��'�8���-+�]= z7R����ɑ?z�}h��n�k�^�u+gHeϳ�J��jL�ρR�&w����}9>���)��9'ǽ�Υ�R��>S���,/��q嶭l����ݭ���f�����
{8��?#����{�d_pŨm��S>V] ������"�J��cb���d��O���ΚAIra�a�E���犉^�.HS���7�+���*�p�;��ʦ�g�Z�j���',�T�K|ީ�|A�2�I�y��OVYV�o"y��X[�IQ���c0%��U2�����N%7M$�����j�9$��Ӳ���J�1I��\� JC*~'p&�"\:2�L=}�l����o�Wxޕc7��+�}j	�����g�W�9z�)�M�c?��.�� 7����.Cw����LO�|�����ܹ�*78�;(��=��;0�I���d�@��d�X���Aꮌ.�.j2�%ŖQOCC�Քr����� ����0�׺,����F�t��'�:�Qa�li��|H=[�v�T�9^F�Y����jH`sV�zye�c���*L�{K���zh�a��y�b�xpHg����ͨ[�{F�,��խ��S��P�X����j.�b :ޕ�φYj�� u[#\���]5�ȑ���n���<�绘��g3z��ң��
i�
�H����^��w.ֻ.��/��G����p �U����$�ϡ�W��`�+SoDdݴ�q�����᫰b�����{�,\���_�>ջ�\�4Wյ���[@Iߡ�2](y��+�kiڴ�:�Z/�?��gW��;��T�6���I�Cl^������X�x����E 7#*Y&�OZ��U[��$��·gd,m��C3�8��:n��hEѠzfh/,+>>Y��c��Gyk���z��q\`5���7]Wt�=L�]��%��@N�!����=� �J����^�Q����صci�����X�xE��m���2��TRt����hK~�S~��UMܯ�]����螺����NWO~8��u�{��o��BX�zf���%�J���6�����_�p�W��#w5.h�}���������j�XtWᄍv���n�ᱵ}��E_��?15��>4��������V�M8JKS������m��O�]TN��C�'��s>��M"�b��������ꌖ�e=7����-��5+4�1��}<f��`��n$�B��l�^�X�PYR�g
�6U���Do��5���W��ڼ�w&�U>� A��~J�g��H���%ʳ(+�l3�ҝ��y.�P���F���2S�sk�����W���J]㓜jL�*���+oM���O&]F?�|ĕ:8d�g�hQV����FU��m�tE{�gB�?ݾ�Jį�Uf���i
��;N�v��̥���YN�x����s�ak��[['��}_��z+z����wu��SD|.��<]p���/��It_,@��̕��l��`&Α��a"O���m�}arj�@7a�����)!Q�]��M�M(*�����k CtE�z'�(v|�]�-�(%b{�U�T�aCA#/���7��+����%�lĸ�ɍ�v��_������.
���^~�f��7��_�����J�(�/�ư����Bw�����2 K��_���bF�F^x���\�({~ȩ��7
��)�66�o���W	7��NU��
��^Z�Fr���e��]Y�^Y����:��F	HWW��Z$Tu�kVV��dn�xG�r�LL�=���K�f9&��䝏p?2;\�d���d�Z,���EiJ�$��+�E���-z�鳍�	=��+����f��;�W���W��j��=��Pe�"�ᔯ�F~R48e$�����*_QO���4j �iG�UΨy�7e�� ��]��d�*F
�C��\.ZY����3���[53W廬�0��8�Α��쵤w�"= �'�Q�n@�h�p���Y,W����G��z�L!ȫ���t.�Ͽ���!�k. :E��U�7_ T�����P��6�ࡤ�b�W~CI���K�������t��X�K<��\54U ��ި�{:;�T��X�,g�d"{!��O���^R#M��}�W�
YN� T��R�4'��2��d<�O8U;Fz��(=Pp���`L7��{K�{���[V��c<��/Z��L�s+{/v�_T)���T�X�Fl�:Y�z��sX��O*�ϼ��
�a/.s�R�@�����X��#�;)��<x���~��qg�"�:W�Ȱ��x���pB����� � 0��>%ӧc��������/�3���X���D^�-T�t��/�t���U���ڵ@��,gzj��W��O�unE��k2:9��(-y��p'�{͆�4J���_�^�Yn���I�vԳ�����Kb�)8�ȗٱ:�f"<+,d��Q���iL8AF֍˾c	x��O}�ʥ���j��K��o�Z�=�s#��]Ȫ�j��ײ?ǻ�o��������S�giy��T��.2lmfze��Q�涚��F+���X�.�*�|��T_G��X2[�n?��U�����F-�'�fz0���=Q ��ͦ�E�R9/���u�~&���2	*���q}���)���ȅ�sx
\ Ns�8vVU��6@��oa�]J邭l��)#�8�$�����.M9Jۅ�IH�o���\~��+/~��Y����ta�j���ҳTn'���8y�d�x�ռ����,uu`t��F��`�R��ZM[gSN*'al�#��]g���rj��ϕqS5~��MK�4;�:�;Px��Ƥ��L��z�L>)�����,���R7Ss}�z��R��͝B˒�6@wP�+��������0N�eb��#dK`�M��I}E��Lvgm����*Yz���?�Y�py�
�{ź�u��/O�*�ܢ>k��+�#�PA�wLyJ@5��,�|KWc5��V�-��{��z�LO�N�Ֆ��T=�{��l�����מ�\Y��K�O4>U�^�V�N����<^�-	,�������K&6�<2�+�zL�1\/jM~��ܩ��0��Y������y�������z�2y�����M�em�6�Z����GU1MK��U�Jx7m���u��3����@���`q�_}�BI
����U+p��Kb�R6rY��^#�v�͞��8`7��7�Կ�.����L�e�ߥ7��땂�n�f�UR��*s��pu?�ω������)����`T�WOS���}?QoөM�X��G�[GE�}o��VP)��RRQD	AZ:�c�!UDA@��D�T��n��y� ���]�Z�Z,�?��s�~���}�9wR�W�,�ˠۛ��&����G�"`�P� �>�Cw����>�[���^36���W����y����F�afRO�i����Xj�3I�o��lu����0��{`ڋ�zj��>�I�͑EN��+���7�&��Iw�Nɉ�B��~�o�|t�-_?戄�v��e��HH��d�e�U_����ӕwB�U�eH\�tU����D%v�0�EH������,��7=g_X}0�n�	[��C�B����S�'�{�2
A0"-h��]v�����m����E�6�Q���p�U��	���a���������r�1�ₖP�l�;�y���1~�bI�b��Z�X+��­~�M���%�t]��iv���v/���?|�ǲ�k��}0}�/����&O '�u�œ�<�l�#�R�G7����y���_Σ_����#�LCi��ܕe1K�Fl�5��3�*��L27���9QZ��+�L�RŁ�>��0�:�5��4��6-I^W2�I��"���+�/�1�%߿���c�G�������!�x���N�f��Q��ؙ��=��/<��b�-!5����.�p0�~p���*-�C��V`��8���`�C����Γ�������z��_�A������.��K���޳�V�w
�A��Vя*���p���2�s�%�6�a�ز�ӡw�~�WÄ�����?*5)�7<1?������d�P���x����dw(��T�� ��,X���$}���~�<�?�q=�7�Ӆ�/�IN��09,�_�?���߁�9�@�A����U�^�Zr�}����E��G1�n���@�'�;�8�o�!�����_ʃD�͋�@V]iߔ:DZ�-͆�v��b� L�8�$K��:j�;�Tȭ�R����9���?muH�
�"~�[��"4���Hq;�82J� p���ڶC���P�$�}k^'���ݓ��<5}"�W��W2��uf�^Uq��|�N��4=�&�gp��h�+Vo��V9�ٵ(�I���+�];�)��?]*���'�_\�Y�<�K[�}w�F���(��A����%�b�3���ʠ$��;�5�"_*A�(���Ε�[q-�%zS�Xe���P�o5}�o�7�crq�;��D���`���)Ef�o�kt�������:T��?���%6j��LP;u�WVB��q��K��9ȭ�Y��\?�J)M���c%�{�],"Pl�M��n,�%V'�z��OTU��_W�V���H�?rH��'
�T8#��3qq5T�{���ͫٞ"d�A�t�����*N�QS�Hc~�n��\���	� ���X=�1��xg}F����(��.��;;�DrXBz�u8@z(0<���̓:y�H���9Kf��>���~���r	h���[�*�~�����(�J��J戛�
��������&94����Nڪ}����Z.:��7x�pd�9:��zX��0dDKz���~C�˚�G��U�GȽo���Q�g�?v�&��[R�}x�����s���̵��c�/�{��������ݚ���1����v��_&"�|���+5I����_�-J��i����2��Ǉp�	V9}xO�5=�X5��pl�}"����|�)p�(f�{cX��/��5_|s����N�-�[�ooa�v:�;!�I{\#[�N�P��LoSm�0@/)/'�I	��Ȥ܏����:�*�Я�j��L}��@cM1��1��S�FK@/��&X@W,�œ#j�{.�"�$�Jɰ#r��omy�/���	+u׆�:ҋ�?��5蔿^S���
fJ���Ͼ��s��*Y�b�b�0m,T�S 5�����N
���@ORG�XO��9i���0���G΂*�7">,����֑v��������@�����r5����}��K���ͨ�?,��[Y�0|*�z��s��u��O�{H�^�e������ �5l"��\,���e-=qa�7��|�]��+����J��XL�0a����R�n���-�C(.2J)�� �7m������>c��g�^�'n�b"׼s�ɚ�c��3��7]P����=ZyȌ{F��/ɧu�S�We@ڝĚ�i52��'�=Q��maQߙ$x�Xo}_yK�dW�v|��o"ν�_���jE��ܠ�Q��GZ���:�pc�,�]����BRJ�I��B謄ui�s��F4�
v�������0z(�4��rқk��"�:A��I ��YI?�-8\��c����YH �27+yL�z�|�h��7��z�rD������_��S#Dɓ=�{�4Y�u��?������*�j����w A���w�
YG������g�¸8_؇��{+��P�w̐3�Iq��k'5��چ�W��CW^�1��rP2CP:�Q��X&:���Q�G�<U~I�_�K���������E�<pzs��S��<a�m6,&������U	������RM1�ֽ8a�8��q8^M�xh�D�CR5�$W~��W���?!��V���fy5*��)�~L�KuSRn�Oؓ����R��H�t~Z=AnW��)��S&i�d�6sk��h���1N�'#Vë��$�54��WƵ���(Т��M#����w�{��Ί�����Q�OO��z������e><���x(�H<0C^nT@�k>}��`�l�@�����V {tKQ �VQ`z�X缦��-ߢ�ҷ����M�>�p���:,HۻF�;y*�1<����B���޽��g"b>Y���0<?Y��{N��"�U��y������O�2M�Gu�V��)�����~}d����:[��7(?	�T��C��R��@�t���ڰ������}��́2�2�|�[_�+��~���5��8$��M謎��Qe�;�q����!��1b��r��O�F(}��}xeܟE�d�y���/QV�$6a�=�����_yxU���ە��bz�.G�tBi���
�W�XݴGߤ[�"`�EB8�~J��k�h�?��ghX�Q��!Ng�3��Nٱ��U.���U~Y�fO���з�:��h�!Xg�5_�1P�LA<�}�˩�!���F/�uL����`�gI���S��X�j�����5ź{ ��HC V�ȓ�ޥ�N�hǥ�h,� ���Y?�Ey�^������ۍ�	���lZ��u��S��zӛ^�8�v��:�_ƽ���@Sb�oNWRA����i|�蕎x�7����W��R2+�]����@����Bɶ���x1k�*�������x�:v���'�Nw{k��j����:���	�R~���K� ����1k0(z�!,D�)��w���<��"�7��J\׊�L~����s��B����@p��I��uL�63�T�h�+�"��h�I*'i���kR�s����xo�a�R`Q|�&���V�)�41��l>5A�yޜw/R:�F�1�S����N�vR�HC��t\��y��VE|[��
|t�����o[���#=�)PKh��,��&F���� �Μ�f��O��(9�'��[Oz�����5'��C3_�d��f��eߝJ%�����Z�Xެ˸�R�����@�x���Q���
0dkS`ޑf���ݾm�S�s��%A^g�c��2�1�meV�"�1�qf�v����j,�f���F�%b��)���8<���HS+CLVoC���_f�Mo�74���T$�ݛUxR����;$w�mx���\v��C��G�3?�v�#3��A. �x)t��_$Z�@3c0 ������9�������4���A'�@���܀dz��}�Y�7�*7��L7Ĩ"�;�e�J��F�:Eg�4�v���S+��Q�T,x��tv+��,��Ӊ��[�f���9\n��Ŗ�����DG��W�0����f��<���O:�F�J�p�$G0�:lM�	�M!��r�JzY��wAῥ���<�ڼ���"~A	��u:�VB*}���m껨�g�	/�Go4��ՉG��E\�?`��wd4V
�C)-���x�0I��K�eB<Ü�#���$��ώ������?_�w3`��Ƕ�(%�&���=K<��������h٫��/vew��_�u�|7���Yb��-�<|�a4�1�)�m�
��/���f�x[������p��
�ı�]������_�y��0�)3Jx���C?6�[��ޑ�q��
����n[Z��8��o��:�	��h����ȏ��K��ֶf,o�W����5J/��ٛ��u�?^���p!�,_-T�@~�N;/pK��>��^���l�BtP��[O1���(�v���,��9����y��9:1r2?=��[�)�'��+uٜ1��e�2C�{la�v�ߟX��Z�y-�YT�󺺇�[x�q�珠=���b����)�a6���j�R���
T��e��C�F5�9�Vw�NQ�ɪ���1.Ƽұ��Y�B<v>����q��S/�(�����}�~c&��;��"�O��� �g�~p�l��X�"y�Jü�^`�w��4�p��M�N���AI~��#s\ڸ"c�m~z����H���"E$e=w{����dQ���Cl��[qm��ݥXI��W�����X�VuI�X�V�u��m[�9�&�e��;W�?&>���h��?��_�*I�78=e>�|���s�	�B�8�9�� 1�g�s�u5�Aѡk���j�#��N	^��.���L�P����c�+�:#�6K,��^ޖڮO��"�"��[���1��Z6�s�0����"��:m'͇�j2�/68b����`�����](�9�#�#s4ڸ�UX'�����ee��qE~�zc��网cP-�����}>ъVn���N�`i41�n���.ԹXW�H�+��0>�O���_Iܵ��k�,�.���9cp�o�׬y�Z��V>]NlexE�
�X�}bW�O-YB���a�-�L�P���V�+�󭎩�!@�����=���U�����*�]`jM����ў
��wu��ĢR�H�j>���ʛ{3�Q��;֦�w�8Jo���:5�ɖ�k+�]�7��9�p��5��ŗyYQ��7�xe���J��*+��T�)�1���U�/G�{:iE�YJ/�3�V����e�5Y��C/a3"�,����%�ߐ3>m�BM�D�wD~��[�IG{��������[Smd~1��E��T�07/&�kS@#}��Ӄ����ra������f�O����i���K�AuÓ5�2�^�V>�����������F-�!�G6g�|������EG��jP�1mPTӞ�&,���y�{���94�Ԡ�jl?����s7�|�v'緈���掃4���9YRj��)��_E1�%���g��eTd65W��~�	W���]���͜窩>�rvg1˖�V��ޭ> @�]�B[]�Z�S3�O}�� -��7�\?��q�'G{4Ѝ ��y���>W��6��#ϧ�J�(��� �`�I��*h!P���ޙJ!��p��;)��Wk>��eЇ��W^�apn�l���D�{�ܜl\���fP_�h��Vsy-j��"X���_�L�Z� �h�9�{=VP��@T�2=�s��}��wz����Hg�������Z���2M�����9~�
��U����4�ߘH*0�'H���0����Y3ܴB1W�!��^�÷��砒�1����e�3ы-��OmS�C8�[�~�p-�Z�RR��wϡ�����rǡ%�G������|Z�=@>�e�����6��ig�0�[�c��RT��fw%���,P>�+����^[7V9�R��UIP`�}�x2�=Vbu\չ�}���*`���Xh�~`m�b,�
z���''.��>oh�;��Wϥf�XpzbR<�������\Z�D ��,��c�����l�3#��y�N�g5�.�y�vqE� XmT�M���9Yb�ƌ�;��h�HJ|E"�y�Z���$b[qr2z�5)�$`���x�wWk%����&���é�9 �0~�/}�(X+��gh#�P5��di�@����5�Oy��8����f����t���Rb�rKcѷ� ����>�hؤ���jȥA��+~U��<*g'Ն��0���*�6��NB�]���.���_,��5��}�� �'z�l_xu�ָ�-MY�������W��PH�h�����>5b?@sf��]����ٗ�i�J=AM�N�S�>n�$ӡ$�R(���ICąs`nwL����*��R�:c/^82�gaA��O��:MqM�eA�.$��J�P����0�K���z���`f�� r��˿d�u��	L��f� ^���a�e�#
�u%��>phYYBGU�&V�
ڢ�n?���u�nP)Ծ�yI��|}���Sy�l�)��8�u�毲/A�O!�Z_��-v�a�FI'�R�fڭ���:D�{>x���������Z3}д���3��wNab�i������_]ޅ-��:[ʮj�c!{��Q�L�A��zs�۷lc��D������Wա��(Ekh�p�Εq������:�� �N}�Ӽ�%GW��ق&��F�J`Z2��Y+s�pu��|�R����\i3�?jD�d%1s�&���O� �7ۨ�m'�U;�ټ���%�4�D���64ّ^�g�e�E���T�����{�L�^�3c��S������'Cb�2����d@���rdC�fx�����e,w�|	��Y���.Io��9Xp<)�lp��wb�r��n�Gl`�e<X��n)����-� 龜ص�w2�_qF����K4�7N�x�� ��b���8��8�C�'���H/�� =�m��k����Ӌ{s�? ��_��S��ヨ՞�í��n��TQZ��:�~�3��>c�=	H_����}o��q��҅*^+ٰ��U�ܱDl�y>��O��g��UlC1�ݱ��e�ZgM�&�H4L�x>�嚛5��ѿ��4�S`�����nl��S*��f�>}��wt��]���36�"#�yO�fsk!!�6ٗ�*��h�=9��[��-���^,7E�������������&�H�z�������,��|tr,2�]kŦ����R��<^���U�!�x@̲I��I�3YQ߬Q��5x�:ܰ�m����^HJΝU�ȘO�# �G);�]|����Z��L���-E[m�v�A��w	��v���EI&�V���^b�1��+)�g3)޷Um�Ӂ-=�E�+>3�.o��B�o-i�޵E!k吵� ż��y^da����~�2��f)���Z����������s�KN�e����w��s �Z�0�X,*(A@�y�����u��&�����)h���<�p���*�`u�,OM�X(�-�{���D8�D��jS#L2I�a��$�?r� ��Ԑv�l�H��;t�ϓ<�����^(l�;D�����@�2���Li�"���L��
*ڡ��~z"�)��b�Ƒ���%G��].P������&a<<kM���}�5cЎ}g�1��*�%6��>q#R�5��)���!�����E$t+i���k�p���7�o�}�*AݻQ'��'�G���K�j���9���Z3[̚I�X<�=�XA�����-�����_>���K�D�S����?��[�*�5s=����&~�IFW
��j�{��p��s�����Q ���Lγ\QrZ������{ Tb�K�y�ɴѡI.,��F�VxdbY%�t'�����]���ED ��1A~��)��QG���ϯ�-*�'��e%vJQ��ԡ�! 
�k�'x����/���š�FQ̒����(���3�@�?{��0���w�����Y���am[y(�8,w�#8�|�:Ȁ&�g�Vv���pr��i��5"�� ��_��P>W���&D���G���:��H:�|�/�4g:�/F)���K�v�����l֜ĭ!T
��W�9�٬�!>O.��|�;���׼Oz��.�d�"��:S�{�g+Tv�@{s�Sĭmoq�*U�\�� %)Gb���^?��e��!,g)��=��¯K�#�5T@P� %]�I��-پ3`3����2�|^��7�a�}��Jܡ�Y���!׀�دL�R���jU��lG��2�����N�F��u�|Ľ�@n|̷>V�y���L_��^Uh��X���j(��:�n}�d{�)��t<���l��H�#�g�z���ţ�V�{�B�/�Gݖ�j�uB���!�r���Xl��~�ֱ��=_ג�8V�,n���?���Xֳ�?MF'���t,�o��'80��-�u�1ԑ����SzF���1��M�2�;E��|�2�5B�2���L$�D��LOh��Wb���N��C!�b((�0>Oy�mH���5��L;���^D��_�����c���h�%���ύ���1h/򺇦���`zc�v�PѦ�{��Y2��C��|d�5e2�� M4h��!�fy3>�Mq���q�֑v�mގe�=��VV;/�sH�rBr����:�$!�Y��~�Z��h�TO(�1���a�wov��x������_����zI�	ڋ,�=-V�v]L�̄�zl(`��Y�C���Rנ��<��0qS�!-����db�r�ҫ�G���
Tc�Zׄ���j}�3�m@����vr�.buK�8� ��@���')�ΉI�C�_83��f�D�يN��|�E�
$T�;ʾ;�z��B��aߙF�R:Y�����F�2)x�|�I;�����kc^qR�$�~4x�ZKj���a�Q�6�����$�����x=���fT�'�����r�p 8�ݞ���X�'�At\|��$��7c��F��`�����lk8���6����U��v�&X��-q�4(k�I_&
�g?�~�W:��e�|��g���1?���^��"���]��9϶�U0>��ؾ���F�@v�k���Ov����^��b�Za�����@�e��ۑ�/��cD��G���%Yc��T#�h+�ͲA���3fƀ�ĉ%�@O2�f�(�U��v��ZL9��n��vNy�Bl@�M��I�ݽ�ޓIIr��3;��3��bD0HS��ط�N��6�(���P{�\������fj+}Le�զY�����k\�����uZ5'z4�<�[R`�o��t5�B����᳭��M�Y�>u$D+�L$�-*rB�G�O�H��	���o�O�#)R�Œ}����]m2Kf����
[�W�j�g�Vn)ۧ�8�\���؍
�(	�A��kٞQ8�  ��zt���%n�RQm^v�݄O��#QBd/��w�K��.�	�e9{��Dz<w�S<�%�_�Ր�	�v���C_�+/A�A��t����/���:NLd��+:���W�<S?NN|����ʄ�}c=��31vS-���[�e,��K֖�V6-��Jgk�b��sF0�x� hΓ��Uo�Ks���n�Bd�Ϲ%:6������W�Dh�Rx+�4X0\^�T<XL�l� u�}��[�,Y�E[r`(��,X:��N_�p���ɳ�a��O��ݻ>��.-����,o���L������Y��=.l�\��>^F}��D�tq�`���%$���ΩPQ��Z��]��E��1�"�7SDi|��UH�|�GY�:P(	�0N���\<�gip��t��b��E-`3��X���g*1G�I[�Ү�9'��E��!�pSX�j����f�h���`��� �������BU�tK�0-��`'{��G*�so03^�E���_�ꆮ��>ڕ�����TP��?q�?�X�JQ��F$a�h�#�Η��.����8F��_��3p����SK�Qʈ��C׭�my K�0I�=V�0��_�� �F�����Y N��Fov����K5����jF�U�m|,���	�pse�Ԩ?�z���Q���h���0����<,�|��=�4��mٳy��SG�����щi �`b�3s4�L�R����:��!k�2���)^D�si�%�]��9?%�u�?�@ �6���o�ke�����gȭ�6��h�?�0E���$E<`��0vy�B��] ��ۇ�M�>�Fh-※�Ia�a�zO�-8�(}���/����#�F�tS��X�)����J)A��y:p:� �1��)F5�7I���
���������g�ptíTE��{h'Í�T�Po����<O��{Y􉂑h�脳�dA���kZk�{��e}VH
|_^-�t�|uR,q>�(4{i�e�/�&�=K�:<�v�܅�U%N$^P��x�S1�F�Q4OvϻϨ!�Ake#��U�b�c���&�3+)�F����e;�s��j�[/ZX���ܵZU]�9żF�����nc�Ջ�'���[�J�g�&�"ZO��ٕV�WfτM�L�Z��uܮ�e_6�U2fqu}��Cz�&���K�hy�r���k�E�		ے5+Lh�MÑ��e��Y =�;�$��Q�?������?��|��49 \�m{V6ʮߨ���~$�%R�o�����o��Y��P���ӕ@����T��zC��f��Ͻ/����5-P��X�dBf~>��u�~w{\�s��P�½Rђ�yQ����IЩG�Y��|�7'����e3Ǟ4Q�T/
�ݚ��F����i �
0�ʣƳ�nqϑσ�d�1�%t��/���7��]��i8�b<�X+k �4z3g��'�Ɍ�E�����Y�Q�$�_]�`����2��꣹��˷�<���b a�mi��Qm'�A�����b��a�Ϗ��w�g��QqXr��T��s_ �����c/ஃ!=�W�ܼ\�"70vy��3���0�g�ٸ$���������d�Sϛ�:��-c�Uf�,���C�:����������|W;I��{�i{�������g�n���$~�/�G�?Eo�������ˮ��tg"@��^JHyEY�]���K�*��\��5����l�}[-�ϖ<l��J\>05�/�\k��-�����؝���䠐Թ�]�s�4�5Ņ�kh;=+¡��^�G��nu��N�D�T��~��~����7�z.�dF�qL&j���R�
��,T���k7�KG#:2@g���}&�z�5�x�U�m�i�	&`�l
����efa������+�]Y��1a�qiIv��^��7��u��$H�¡�xʁ7�;�8)E�V�E+������T�i�^�
βŻ^�&K�b&ׅ,r�$U_�`=�Q\�S��=KM�>6��h�EnB_����{ұ��W�uԡ��~��\��d�u%�Fz�v��v�HU���?�`��Y������ƁQP��F�������S��W��#qe����\/�����D}n�����*�37d7�ʕ�x�uj����ݤ|�P���O�ub_���[Q���r�n��Õ���]B��jH�;ގ>ߪ�L6�y��i}��s����f�G�Y��{���6�'�T�q��çvo ~��\:;y����cqEd��f�bz�B�p1��U���{Y�}YZ,)�M�H�y�7�cRo���sD�q��"��z�q�x�� ���?����h�V��{�]4���D*��G��������) ��e�Ϋ	�ل*ɒ����ؿ+Y�*L1�H�/�Q�O�9�_�@{U���1�޳\��&�����a����}0���� `������4�LX��#<E��EK{he��(-�S2Wj��B���[��>�#l���ߔJVB��ׅ]V�)�FD4j���ጾ���T��^��kw$d���4�:���_��	�83�4�5B<Z�up����,���1�9LQ(r�^MV�WY�)P�j���>b��;d�[���T65�� 2JV�K�3���8<��H]>���r�1/ ?n�O�ر.�����Nzt����R���O����W�Pn3S����m��]]���w�&��?���3*������%�5@��ñ�Pe�%���a���Z�5���� "��O����5C�E�B_a ��-rZ'��zMuH*Ƶ�=+�:K����j�y��g�o+��у=����iB��I�a@s����hϏ��Ƥ4��v<Ky��Θwۻ꧓��z�Fp����|Y>"������zn-Y���WIw��+�c�g\ _Ť�rLY�k{���8�B�����������d�z�Kc?�$��[R(Z��9R=zz��Bww6�B^l�\�!��U�� �;�y�O��w˛�?��<H�e�W�v8�K��BZ�A�wtf�;�@eem�����_�O9�.}01�*
�RÌ�,Wj�sJ�YJ��К���)��]L�~��]=�����w�}���Ώ�O�FW�}-���L�����\rpH�2��ր��+�O&����y7zC��> +ȃ���g�&��V�HV{������p�'yU'Q}�k�t�r?�}T7|[&���P��$�$��>L�'�<��
�(_��߯�S��KS_z)�ȇ�GP%FOߴ"�PF ��_�H3l�K��[�I��p{�%�n��.2��p�����١8� �t��E����c��"��ú(�mhW���--�TԎB�@j�����0�W1	�����x�:���n�-� 1�U͡��!�iYЮ$���ڱM0���X�����h=�
@�~�{�jf3}�w]"1��j�((��D�~#n^�R�|Oڠ�=C��9���Qꌕ0��+"�z����'3sd}��Xb���?����I9�u0[̸z ����d�����������өP�i��ux��R�a��O�[��
�񾺖�w*�z�
�?%v�qL�Ƕ�DP������B�,i��E���>����k�Y"q����?Kó4���E��5��I^�8���^��.2��ho<���ʞ|�Q�r8�hem�7M�zͬ��zl	u�������M�ǳ�u�d+V1���"*��ec�p$�����d8�348eyH��J����J5<ֽ�jrk����<�Ӓ�	��U[�t���M���Tߺɖ��A���k���(2�p(<�	@�ee��I�M+�����(���_F�,���0�p84з�R�e�t��)6a��3|yK�y�o�J����b��#����,����@�?�k�2lО�_�O���-��w�բ��u��$.-��⾓&a�o>C�/���>0��p�o� +*i�F��ҍ�"�0��B�~m��i���+*�#n<uc��&��ߗ�楒����//�A�wXR0��w��c܄��=�Q͇
�A�����A��w�XcX���+������������V<�n�t���7 ����X����s2=���BK�,y����h�l�0�sզW�����C��Ä���/�t�R��+0g��lar�gկ��eiӽ����O�q�mk���v�<�<�%�<�hy*-�}Mk��!�V��0�!��ֻ������k� A�eM����<�?�!�>3��Gg�.��X�&Pr���l�'l#U"vt�Ɍ���^(]�N�`)�����oJ_ѝ�����`�Bn��{�9j��c��T24x��L���-FX3R<���^�C_������0�Ӕ[���9�f�Gy�78�2��7�k!4�Z��酆�Gi�Ҝ�e?��/� ���޽����`��y�(-����h�ٟ)�L<��0��]�8]��f��U@�J��˦�~�d���o��ԟa��)T ���}a�w-��3���F��L�A��]�yo�Q~Cl���Y#��x��S��h�\%�ً;+r:,d4�*
X�tM�
�tP�Қ�\)�
��d��l���Ʀ���/k@a�<���p<_�l�NV�l�B[�
%J�����
�x�tz��n�o4�`��FϚX�)ZʶO�34֮��
=�~�e��t��r�u?.Epܣ�خ�P���U��Q��<�N���;w�\�ą��a������A�~�������NaTW���T��p�샳Ǡ�a��6�/�gI?(yf�yOV�ZD}����Cy��ݜ�I�����5n����e(����*V��ѹRɐ��2�rFg�s��ߤ?q)�	g�;���0�2a��&'�g>>�ٯ��S������C����(�;��=�ҡ����~./]�r/�'td(���^~�y�a��$6���!'���(x��n�8נ�������m���8␝"kje��Q�z�$���UR8��L?���}U;u�f�|��'�	5��,>ڒFy�L�{��hIJGu%E�06t	/Y'0�]���ݻ���D?Q�Lhu���=�g�8����<��ey4�3���B*����	��d.�[��������66l+��������-D��j�}���h;��X^��3㽹�#c$6����͔��U��<��~쵘~��ߤ��C���q�q��q
�l{�%l#�������猻�R؁�ԩb��~F�¨�A_@֯JOK�6"AZ�m���'�q��u�Ou��Z��?^�>�l�=(6���Ƚ��S�#/���F-�qȚ˰��/� ��w�,��{~�,�Z;�!�����(s�K�pv��� �?wI�A(n�1��8�M��d��\���P����v�W�G���0ه���jyz���fF{�I�M�dB�p�/�����"+2.��L�ͳ������{#����t�φ!<�cl�w�T0��X���h~��-��n\1nM �t�]p�~ YTgs�F�1�b�'������h�J�<za �0}�� �-dru}��e(Mw$l��M��F�:��$�|���qQ(�`�v�Fӏ�'L�O�ʣ�����p����mh)��ign��<�7��٫ҌF�Z_�4"Lb�,��
C�����u����3��9:t�Z�BP��h���Õ�2	�=h�Y^F�R��5�޲�	�ݫ�l�<���Mҥʻ���|�O��cK�!���sUe�T�_@w��
�H��G7c��V;r�7GЇ�PH����(��T�
��E#��"��7/4P)"��;E��q\H��z��K�e��u(���ti����Y��b��?�ɸ�c4g��\��o�ބ���L�n[4�<l���(=J��B��Z#���	��>�<[V���QY��9e�x\_�h
�_�8�ФzO�{�\>&k\7�ǥ�8/�FK�=:.�%�?0l����=N�/|��s�,��F���kZ���拫-���1�Ay��Y��ppT��G{��)ǭ�2O��w���'$�����D��u0�Ro��F���`���5{G�c���}�|�F��s"C��S���	#גs�R��Y��	9E䲲--��������38a�&����;�e �#���L݀�� ��j��n1�g�s~(`�
���L�>,��ѷ��E�'G��}��!��!`��;'o���_��]λ����Z嗵�5@��ſκ���.�NGLt�g��ͼT�`iݍ�=��xٚK�T�-�	d$�Rv��������`�W�J�����+R�~N��o�]n�<Z���g�����x����@�r�fe���̉I	ј�it�Y6���Y6_cOy��`��Q�����1�f���ᎏq/(��$1P>vc���O�����C��p�.Ӱ4���Pŀ ����"�#�in���F<�ү<����H�m�����}\�������
߅�H��Wq��kx�N�3O�t�i��6<��7���r���/O� ��5H����D������vS��M�Iq�y��P���l�9d�����p���,)�Xޤ�ﱡ�s��c<�I�Po)]Pk���
L�J��{�^t�y7*Yv�#u/��(��_|U�N!%�)KJ� ��g�UZ�{A�j��M12�_�8%�?f
��ԗ8S&c�D�i�@�*�Z��M��V�b��_'�7S����PY�3ӛ0�ú�I�;m���!�f
e��S���#�x5��%�~��P ��� +>&�oX�\_M�L4��{
	ޒ�Eܲ��� -���sV��V����N��j�g������[��X��s^���o���ը���{sw� �<��(ǉ<F5;" `c)V��`a-��pZ	C�fyWD=@װ���� U��9�&�x�OR�|��*�!~틄�s/�Ү���4�g3�
��9-ұ�F�-����h�B�v]�g�)�v��Ȫ���3���}��)�L�h�L��K��_g�{'�8w�{��q�}hR�?���Y�H�����VC����+M���I�vߡ;�ɭ�2l����|�rХ�|6T�J	���2�!i��w��������b�pqC�BU�2q�x�/����~2��N��Ca�3����S}�� q��{��,�����0f��B+1��Q�<��*�N f��1�U�yj��>���sl$z�@�*������i�h5�}��m��<�x�/u��h���)t��9����
�t���b���d�3EF9$S���c�ISxR4E�pH9n�����2ʑ��8r�PK\�����<�aխ[�E�9��� -|�1�&J��p_C5Lԟwh�ݙ�X����i���8axS^��k��]���`c#�Fp����'�VΈ&���>��b O������㱝��OdƎk�[l�����q��O���?駶�k��`�#H����p�o�������-�S��HDa�`=��S�����]�zw��l��;�p�JL���,Lwr�(���X������LЍ��O���3��ih�t��%BM���L����{"�ຍ�z
�~��OKʊ|5���+��Z��}��[�b������^�zz8��WREF=ػi�`}�q|]�|�����"�w�cO��E�o@�����7�c�S��}�73���_F0q����.�(��ge�}^�U�+|�Jn�v��rZ��!8ꟹ�Da�ގ��p�ΪD���;�I<������1�"��v�T�L���qM��.J����x���:<����^M�]�q���QaT�� �HA�n�HWi�T�5���
"MzJ�JP)�Ez�$@�B�=�2����޵d-��$'���{�'�	M�_XM(1>�� =T:�{3��m3������$���G�v������2E�����0c�-�[�C#�rӅ�R�_�[���/��I5٪�x!�d�&�Ύ)ah��M ;H�ޑ���Sۡ���/-\����߈�9�R�p}-R�1P2�[��%u�p�C�#�D��J~��B+��VMf�(�H��s|{0����/�.�m2W��3#f^H=?=qH0o<Ua��L��[������⻌��*�f}��<h��.����$n�M��5��T�QL��]�����}p��և�K<Z�ɼ�&��]�J�اT����^7���qz7Π��\]R�C��D�#K���p��I{���2H��<BG	߃��á)�:�����aIó��j���|�zh��ղ��R�v#���4��o���|�9��'�.�d�`�a��D�h�۩)�������[6�ߖ��}Ѯ�^�%]+�� �+O���=�����o�X��v��?|�ƪ�)�����!���S!�oFo+��&]u5_$>�׷�}ߓ��`o����i�^d��4y{ڜS��y�
$����G���ѓ&�C�Bg�3
e9�el�L�:_l��>����^�5�?��q��f� ��$�_a�ߞ��n�5)��~c�>�Ѫ'��U��J����ѥ;q􊐎;5vhR�J�by	�N�4(\X���`��I;�I�]@܂%Md���T�3�2jE�ij2����/��pV����!v)�O%"��eRA�É��e�iu0F���HW�U��M�7|Kܩ�G*���+�����5�����^:{	0NY�qC&
?qyo|���׈GWb�iAsz��=����臙�����T���F�i5�W!�y�mr�> ᤿sa�g�M�me�&��V���N�I��y���W�%�zG������?E3_k�ܙ�J-%�Җ[��[{��Y0T�E�2�3P�┌U�i�C�9�|, �;��_�n&}G��S|��`�w�i���p3ǭ)T7R��MUuB߃���c��6E�?H������B������_�x[h
�Ȑ)I�Ǩ
P��U��xz��s*|��ы���m:#>���/>���T���}5*ݧN�L\��|�C���%�0��))*/w�Yt����#���B��B�2�=u�G�v��T,�0�D����?bN�?��O�CG޸'?>
�˭�жh$[�Y�4:Zr�B��_`�EDi׹���ѝ����/_Np�LŊJ�M�h;�]�������o�Ve��6������H�'Ӿ�B�#����[zw��4�j|��У�� V�F�P`�H��R�i���s��lg�ZM6�0D5��Yp�0l�rv�咫z�0�E��W�?�Ƴ�V���8{\��n<歅u�.�<�]]w�H�)\�"���@U�?���!��x*1e34�K��V�R�z�-P�j��������Z�g�܇��}���52|P�3[Vj���G;6���h��[��{�-%%m���ΓIߕ?ԃ�fr�Bj�]���C��-���@��e��j���4d����b��߆RGK�_l�}��٠YN��^6����؍��I��'����������{.�F�g�3/��{;\��Ү�C��(�x+���N3��z�;��e� �x��^� �T�k5�~"b�D]i�'W�&�y�c��5��ª�O��[wbǆ��0+�kꝄ�F*"
,�W1ˠ�NxX��v��0��:*4#�UU1F~��<ǂh7=�A�zh1%"��3;���ݦ��i�#���W23���3�oy���d�f
��և
�E�F�
�/�/P��Q�����Ƀ(jBQ~�̔�`����h��f�2�gx�O\�s��Ja��RK��򊳒��	01Qѡ#�#u`b*db�+�_ͨ�t������C�
�H@fu�B����eYv�*s��kNn�t]������G(���%e�	���[owE��6R������R�`gz�9���ֹ�w8	Ɂoi�+�����?�#�p$H]w� s�{o:@-,�W V��W?��SF6��5c99���	���C2�	�@�>���2u5ժ�ϼɲ��8^�W�݈�On��=46TZ�Dg9)�Ε�Ӑ���#M���Z(���`5lTK˟���m������s�)�<��y#��.�:q�':kD'�ų�%�=p�:�B:]���������?�V���5�	4O�9W�a7�ﹹ9�e _���ɂ�����W���J��t˄8��b��n�=_���g4�yMK�W���DdZ�]��Qnntr�����A�T��f��	
�>��3Tga�hܷ
��o˴Z�� ���@�k���Ew�}|Z����l)��FJ��7H]�o�`�/�]zM���([zJ���d�����1\�E���7�H��DB�h���ϫ��{�֩ސ}�
����M	����Ѣ|�Й3h��NF��؛���YW���ɯg5���썢��
���V�Ţ|� |!�o�K��ؾL��ה�}�ᢵ_&�������dR��)��Y�h` ��f,�	w_t �T�J�PT�T&�b�I�g�X�,<����_+쌨�R(�5?a���o@v��
��u���r]�bG4���G"=F�]K[��28^r�k�X�V�bۭ��2���^�@��#�(J�eڀ%5��[�륍.ҩ��l^�!k_/[�^*Ȫ���x�1�݇��9�����?�!���20�͗�\�V�\�'m��WIώd�KS�I�uN?�x��u2�aXf[�FY�`���'�8ot,^BL��xɿ���\#~�K���n�Vj�E�!g��Ɠ�L�j�S�^E�^y������~k�.(C�y)���.��A">��ލ�(��,�3P�}�v���o@��W]��U9���ۦ�Uf�I�0[W�:--��W�9�g�>��!a(�<~���xR.K��M����2������ʇ�G}5���;����C{Z�~�G����t��%ԋ�
��rzߍ�t2�
��Q b��<�t��.ˍFD?�}�gzW�����٥��f��f^D��9R�:I���Jo�4h�n��'�S�,�����1�� ���$g�-��w"��`'Ҥ�ٸݝC�{�IUS=�\H�P.,4v���$�EE� �{�4E�������I�pL�����h��5��@?A�֋��xx�І�s���J������+!�o�t�K`+١ӣ�^t:�%$�3����^��z��Nwy3|:f�\Y�2�Yh�y2a�f؁�y���-Y��VJ��J�-����X}���EN]�g�[�7��K�>R������� ��Run��m�E�+�uN���7�	�24�zM�{Jڅ�<s�0Ev�-�V(G�4�t��`���n7K��HN=8^�S�ZE*����"��̕��}��N�O�A+B:֌nC�/�A	��������h_�Bgcц�E-͙�hkG*#/Ln�t=(��Q//:PnTN��S4���$Y��L1���y�.�0�_���X
ʞ��H�/��'�����v=�H���p|q�GP��jD��Z=��Ym;t���`~;��qH��z�ߗ-!?�Z1�0bS��2�J��v��9��>�P~�#�0�6�&�#��4jav��Yg�!k�7���$�t�Zy����羫��t�0!���M?�7���*��h����A����L|-�3&)�z���!Ǹ���֮�fC��AA�^A!,Y<В�"�R[h�6�M�� ���{�$�9cCy�f�߈�<x`ad�ꏞ���>f}e�;9��0�e<2�~w���K�>�V��L0�dC{u%�4���FU:2/����S��-�-*�i�]��<�u��[J���#Lj���aX���9q�(�
���`|�P�����ށ�ε�J���(I�e��Vg�ԞS9�x>�h�L�,3�u�|.�'�-'�vE�Á��<\uCU��<���%E8�4։��k9V4�,�3�.C��&�����Bڝ�S}���}�f���V�w/_^����q|��~�����Vm�o����8�Dp�z�o�x�:4u=umبb�߮Wq�� Uf#&�a9o۶�/��^JD�*;�ӽ���̈́ݰ�4�;�z�g��@@�;��"z�w�HK�@9����Ex�~9f��R.b�ژ'������ca����f���u�wN�BF����J|�J�w��M�+��#�Bh��/�4_��mESa�G� �_RT��T�"��&�e��|���F�I�����N����902S���[ƣ\��x� 2*��\�|�	/���n,�lkʰ;�S��e!=�m+��e떚��%���N�1�]����2@m��P����Ҩu�Y*�h����e^\��vL���r�b�Z�CA��j����{�/��7��4}Yar� GzASg�c3��^�Ϣ����Iq���
M����]�~90�4K<�yT�����4��nz���d��I��	���\���I�uӘ�߁���g��	3O\^�g֪�T��RB
�c:�A���`+`~��.�WɆ>���=pO�Z��k�gM�)0۸T
�WB�Hx��ݗ�1���M��AH˰!�xM{���]|o�*��Te��O����IlG�R��f	�l���)`̞k������KxY��SI���6��@~M��e��� �	�z㩘������7�_��1U��g ���8P�{IӽQh��.��%W=����A's�d`��_^�$�ἴ1��*�@�>Ogj��l��� ��yx�r�E5�z��3�����3.����������l�R�������4�m�n�{��tw�R��hb�i)�1-3/���(�H��λ��q�������U=�m���p�s�3���f;+[�_��qH��� n��q�:���e@��쎺 )GUj�՗tq���%>H��f9H�R��:7�����̌tNT�=�9���aer�IϿ�����Y>� �����o��@�4i.8/<�/�N%|�4����k�*�d!��[���\��d�V�>��~_MZ�i��{K�=��;9CD]�V]��M�|��N���,��`��9�\��rF��lk��
��BL��� #o����nW2D#v���#��Lm���Qf�ќt��qP��X��K\kQ� ��f�h�g8�|�@�]�W���v�q���|r�"��f烒
43�JGZ��َA�>�J��N�>oqWih�+s��Q���`uY��xg�(љE�� ��3l*f�9j�=G�J�w����66Yij�a�t���zs�dcl��;%���d��c':�G"�M��:(y�������͍/~�x�8f[SI@�[�8��دr��3O��Κ<0T��,�Gq7�)=�;�  ܩ`�V�X3��(իK
%��0f��2ᬾS�oP��>��^ܑ�U4,�	-ዼ�-��r�u]����b[[G/��6�b�E��MA�K$m�O؄�lc��)	�?J���X皀�BAO��E��o��;����b�Ө(ic�hW�3��u�_��4������<����w�Za�9C�}<��1COo��W�uZ�C_������cF?=�Z;OˤMwH`���EL1ui�"|Q M�Nк�Υr�i����S�C�A� 	�{o3�ݺ��bl����E�F��p~��h+��=���0��i&,�S37���X��mEN0���M:�b2�28@���� �չ���M!9�7��ϕ.W�;��#,-��et� ������h��\��يv��@H3�������ϱ�f.2��"3����)e�[W��D�H�`�<�e0���JDE^��`9ϱ�Jt$#%� �~��q��`�6&���=�k�V&G�tf�b� -�o�[Y@[�_^�}l�C�
i�-��}���X��g���gm�.�K m��l��]#k�W�.@�A�|�N������`��s>c��N�>�G��oF����@�� ��3٢�R�&E
b#?�[��[����� h,��f5G���� �9��y����9��b�SG���B�۸J1��Ui'�(׼=�ӥpn���r�Μ{M�y ����1��}�����4**bx8�*����%`��~hb`�Xz�� >^C��� ?����n^��@��~ ��ϭ���|�ix�~�����є�L�+Bjxa�b`ty�I�����萺�)yp5͋�����Z��̱k����_��}�T�'���5�3,ɤ���/I<c��|4��V�ݿ�ecK[ӈ����@�Te���L)�$)Zz;��D�:r���u)�ݾD�1�2)���}+��Dɴ e��{Q��e_�|m�̦|Nx8�U�r�B�5'E���˵��뎣0ѐ�o�Ѧ�#��p��m�vG���I���?MF� k��~��0���\s��4� �:"�-��i00� ������ ��vb^�����������(qW@�O�!��쪁v��m9\��S�]��e����0j�.�\ߤ�����֕� �zp</+�������$1�`���q�ps����+o��Z��߀	�c��@9#'c�8���i\ۮ 捾+$�P�-�Y��p~�E
�ݮ��mE�}�Z���.���J�ɀ�{IY���G&'������>{̕��@�{��P�Ց8����0[���0�C5��A�nd�Em����J�3ٞΧ�Hefui�)��K�˕� 򃛉�!���ݎ������88$��$P�������v�i(��$�r�(tE�d	�_��F�\����Phow.e)4�
���+����.����լ�2uvI�]F-' ]�����0��&�r�y'#������� E_��b����Ũ���� �� �ؠ[�����}�Ϙ�J�ĳ����]X���Į]%�@%=��w6�ץ�B~�Ěf6m�O�!�1��G"w�2���( �Q�6j�{���F�\ls|� K=�~f��T�s�;��27�(�uQm� ��l�]����}��q�@�h���\�$E�%�L�5G��)�&"��W���,l�5���pSz�(�252�@��]+�ny�!�Q��{֫�B�Xs��Ԗ�,��x[�x�hIk9�'0V��̬H�I[�&�I��.22g}
�ccL��M��l�/[a�0C�H��̎�}[W�����;-/��^�y��h�mM��$&�! #o�H���w��5�J����X_����!��ii�Lo4���¾<S���A��z:|�i�M3lz��49v�TL�J��{˝Q���?fS�b��Lإ��Q�h<���6�W��h�R<�+�%�\
ۉ�|5p�o����Ӈ7n���NsԨ6?؅z3N�J���<0�+���wVC����҇�©u%9Qs8׿�!I@�twl����5�Ԛ@����6���?��x�Ixcɓ)��n�Ɂ�����@���3h%���(^,�VL������x�UHl��PBkBƑ��a�sb�OM�P�5H�8=ݩ|Ҹ��R1V��\�S��6�Y����hP-�tѢ9|���X��I���C
4��I⯗	y�莩,��$���ߪ�&s�7�=�!OL��ݠ�v�S�Y�ň�.�f)��EL��,N�3��u���gij�����+�ʎp��yd�QU8�+��=����<��H�f'���@��6ZdT�^t¾z9P_RH�[*\�+CA]��9�>����x\jfwy%p����eͣy�UYam>���r'L|����Կ�,�d��7��d� ��X�G��;����t�V`'�����i��ȉ�Rb㘬ѫwo��!��h�wmT����R�$�@�+�6�������MŅ�؁3x���/����6SA��;vu����F)�p�Hb<�r��0�O~�S�d�U���H����J����{3�TfZ�i�
(l�Bv^w��2m�yۏ���� :׊�h�����d��bYLgju��k�6֜����G�U��L;:�W�M��}�*��FMlP�4*��U��eD��Ao��^��Vڱ��?�&?����!�����i����̙^�rY7d1$u���h�J	T��@-0�jn)�۪;�����V	�s�s )^?|+�h���N���W�Q�ٻ`�v�H��N�`T^�����v�i.�ÓJ��E�"~`:L�0��:��n�@��a&6�p�s�u��ڠ7�j�a��[��bGٺ�9���� ܈8���E�e����q�k��{�B�o P}�׾QgEN=c�"\⡺(��(3�V�b=���[�|+�8{p�h���m���*m�N��0w��0�UL=��f�^ی�9����!�9/9��m�'�[�p��u@���{]w�Uo���9��8�}��1�r��K�?�z�N�0b)��B+�z�M~����3k�{�z���tg��gŅT���T����L��HX�]���Đ�NJ0�<��Ɣ6��j4�	�ȋS���?�^��[.�]�g���� \�P%XX���V�	6�E0`pP��`���#�j
�L��4���x�Z���lgB�,9[l��w�f#xN��`LI��s��9�ڽ��'�C�����1d��y�m)gXr���ǫ.�I1���-��.�=�	���4�-E���:�+�,�<�V��Kq^�-��|��)~���=>E��~��P�.������M]�$�qd��ӯ�O�!w�_����E�"z������,���L��ϣ"h��w�J��ï��D)�dJ����e��uo|[<v֛>��0J�#���k�?dC�T��%wB��C/G1i�=w��3�d�;[�p��I���U78D�]�[�,�t��k���*M������ Fgef���c�1'�^]�����u����7��;w�˹�� ���'����BOy�������p���	�%)�w2�<t�#g*6�+�h�?>{냯ϸ�1�m��f�i�@cë���E������0v�6(ɔ�l4>U:Q���{�H���|!%Ui�����ks���n��4�_�L��'-�����B�QO�eۼEA��*kk�/<���yϽ�
�P\�
fm�yϋSr+�e%�z�rJ!���u�O2��QUP����{+��5x�-]�����~�'h`�2E�5T>��HX���Jq��3Tc@f}�\R���6�̒��`�E���J�`�w żyvA��H�\(.��zF��S\{����� ���fx߷��G���%�x�+�V�D�v��MX�� !y�2�$j��rr�[ )��SR�����6�2g��vC���[����B�+��]��C�'��:�����;��S��7� E�x+�oP��R�ߎjw_�Tќ����8��K�x+;J�r���lv�}_��!t�
6l����3Q�@"�v�Q�@���U�E��{<vr�˒���`?��/���_�m��`Ñ�FG���OIh����D�_ ��gP����[�<�4׽���^�]Ҹ	�žbd�:G�^z�m-m�.���������Ƣ|����%#r�ZCPq�	�X�@��Ѡ�������K���1v.�����!p��S)@�^w�����H��O6x����J�V���70�l)�R�[����cP� ư�,��&n����>�,܆���3�:O>����G�W��.5���(ے �,r�v�
NX�a�QZE|q�W��?�.Zڇnl���l�O�\e��SSe7� /�zGb���[�8��8�a)��	 �A��/�*N^�]}��zOiw!�<�W����$�#��|��]ï���'d���s�dN�Q4�v Wj��*yMM'<5\�6a� E�Gq���0���Ygl��<�©w�Z�°,�\.�BQ&������S�����5���7�/5h"��S�drO�=������7Վ=�z?yc�p,D�_õ~%�H�)�ͺ��U���B3� ��ƻ�^�P���{�P�Z����Rg}c��j"^�Op[%M-��L�v⮻�^+j�7.S�9Q�����}��ݏ�څĦ�.��@�e��g������I��VHг���Ȋ��rk����.�ԟ��b�jDN�ښ�3���X�?�&w���g�Db�Q��Lt�ju�2F������M���"����Ӛٻ	��@v�Al�2�"���7�+�*0Nq�=��-�f2�b�`���ޜ6H����
���'��]�u��O����\t��?YE!c.E�lIH�OM�{��X��Q!���%�p���l���ZS
���ۀF�9�WtlS̴�^��lL%)gp�kU����u���(�x���fYE��k��T�����l�A��r"���*~�'Csz}�)�<48g�ĥ�E!��g��E��e�����f�<�6�Vgژ�L��I���c�K�:W�YV���n�uo�������.���i,]�'��	�>ϥ����&��>0���"�b+Pp9=wt�F�`����-�k*��wQ��S+"sW?��ɥ���V�'yAqƊI��lM�,2���l����h�c���ʧ��p)�Ť��~��~�d��w`����)Ƴ������)~���5N?h6����o�Z=�a�WY��k����,��5�˰��ɑ�����gI=�vB];��<EARb��ō`��1�٭��
Y猨�-U�D��>��̜m� �M��ܾ<�r��J�����Bv4"��� �$���
a_A�̦̳S�L���HA��k�f�%�h���yn�T���G����^�chc��I0��SLc��6	��i�wz=�Zơ#��&-9JR��:@�V;��S$�?�0J1�0՞�u�i��WO�߇�E����hKjд�&w��e%Bf}����j�Sm[oyl#V�{�	�#�Q�;}��VC����I���<i	T�E%e��f[�����傑�J��(�U���)|ޘ
��{ "���n\����[�����!+a�b�:����RH2ä��7�]�� ��DX�V�&��Ɣ�:��e2�9���!��ȿ2��&y)v`D?�4�Z*��\ccm��B^@��x��!0�����я1BڌX���Ff�<Z�CcQ���gu�沬	���\uB������p�칑�����)�W�^�����W
�i�VO���U�ec�ٝI=��C��X��1Қ�G���J'a1����ŵ��A<~�$<L�ř��r�c����_�����t��QR�S֋���2-踹gaI�EH��&d�����l+���	߮���a��x���ͅ�๿�~:�G��_G�Ck.ZA_H�~��@��x��G�QY�Q<:L��΢�<�)�~�T�!ݼTu���:i�3���R�@�6�@�k)融�iX���ik���V0��=?,5в2\��Êc�הbV�H�=���zb�ϭm�A�奢��b��������8g�Ҹ�����)`=ᔢ&�Y��EM�w�6W�`i#�K��<�l��|�0.�����1>�	���J"��kTs��[p}�Z��T�B>n��}�.A�M�E��?!�4�)�H�^pߠ��d�N�H���H6�VM���#�gP����.E���ڝ�]ħ>E�u@�m��pX7D !n��3S�Z\#Ӹ+" *L�����s��\/VR��x� ��"�R�C����C%7@������gt��ʜ��Y�/�͟�%�����:I������ǀK#��&$�]����"�m{/Oas���Q��7!�l~�lKYԁ�_oOތt-�&dY�!و���L�^��8q6�Ǔ�+�/�1�V�FF$�������y^����:���E˚�[@k��� ��7�1 �r<�0�jl��AYqr���f�L�sP���UJɋ�R�)0G%I����3+�f0��� ִPI,2?x���O7�Ht�"ĬgQw�ND�n̖�O���1�X`���l���y�d�Im�)K3Ӷ�
1C����Ff�@Z���v����
Xyh��C5"S-���d����7�p�h�릵��C���Ӷ��`�u�B�r5-�Xͥ7��xN,1�Aӛk������o�5��j
w�E��nW�|f�:�$��%�C D+gF�ӻ�S�,�3��B��?0 ,����.�as�چ-���
9������.��d.�`�yBb�,����䳌B��z������Ŋ���FF�?��5&�N�Z�Ī;��EC���p&� !���D��IGM0��u�[�h!�q\��̀�T���[
�Y��W�܏ XZZzK'e~�jW���E��5i��j�Y����@
()&D���G�E����iӛ����BI���r@�j?KKԷ�k�Rz@vC�-�Ƶ�	��ǧk��Voy� �����y�� &8I"�qk�ύ�����z�q1!Lo�l[��l�'jƚԘJV|5�*ԙ�ؽ�䆱K��4��q3Ԑ�G�Ǳ��f�x�����F;�E��t�6.�u_PS܋rwe�c��rq�-���¼�����ߥ��:��&S��e���%ʴmt��X)6^�7�5q���S*�BW`��;2;7������ ��K���I�9����<��YKZM6�N(�$�l��-����G�d�Hvu��+a���(�G&u�9��^,B2��i�rM�JЅ_͋T�����5%K��D�����NH��{)DN<JY�J��� �]���$�Ku��vsa� �m���J��|Mdw��'v���u���iW����4�g������䞂�����l)݈k�I��pcC�6���&T�k�hWEV/�,�4���Ո(�Mm���~���\z�L�i_*%[�:�!����a�pg)�y/`�@���	�8~�&0�QiR�G�_$F-�xIFh2�����/��nY�x�Y'ֆe�_��������h���k�=�Ƒ���\����;���N�Bo`m��D�F���	<t�ݚ�5U�]${��m����kl0v;��v�O͸MΩ	�j��D���&�O����!�S�l��Y�Ԗ�q|�%���˄��VAw�KY<f2=9z�~n����z	!�"l����m�QQ��ޠ�+4ù.���_�L�Gٯ;�E4�;�`�9''A�"�$ݿ%[Ppi�QXx�s�U��	+˜S�GBr⺚��;��-Z�m��֊A�}���`���'���a��~]q6���Y�VRzI�b�&L�#g�K�� ��u˵�C�d�Ǥ?�ZK�mR�H7��Z\M��%�śQ?�H*�yJ�a��"&!"�g,�Z�ӓz2�g�������&3���GN���n�7�.�P��v%{�A���/u�kU���y9�� 76}>x�����	��]��v�ô�m�Ȇ,�ֶ5��6����fu����Gt�\ϋN%�B��b���{�j��ݼ_(,�)6����]�&��bp�},߅�N���#ؐ��������c����qQ+8���a��PŃ�s��؋��1ѩܤ,�Ȗ?A��#z����\�
�.[sg�Buv�������D˿},����c�5��f��1{M�0Y]`X�X1ݪ��*Ks�Bڧ�UD�/<�miHh#��*�T",��fjz��(4�70�|���TE�D�����m��h�}����F�,FcE%����F�/r� �e�Nd�h��0ę6�J���L�7���}��=�Cs*��,�C�F���G<��m�xh��%CE�|J`C�Uu���{�M���Q�m$?H������RSMp:--�3�b�¹A=7O}���'����������u��.
�,
]͵�'�̿{
�l_Q�b���f<TZ��4�y�]�F&���Ĵ�<eAQ��p�S2����r�k��q3�*��3[t���93ٗܖaxu}�y�$��>�c�y��ٍm��c(�^rxXC�ޛv�ʛP��k�`�0㚑�M(�Ƌ�����+�"�೵ZT^a8�쬏3l�x����aYb�*�����=���FD���"sB]��z��p�|�L+c���W�<��@GyJ�ڎe������OU��&QNƤ�Z>*��'����lp��ڃ�ԫ�(�LN2�g����L����_u���/������V[tbs-�����8tS&���&ͼ!����s���P�Q�i����������sǏZ�N����mep������m��͙,�K��﹪��($�2���^�}�ìbc����ɨ��\���G�e.�b�M��FZ�Sf�r������>��S�0ӯ";��M�v��ڀ#���#��;A)�/��6�]'�D����!�Qwv�����mYzn+Gs̝�J�u�,,Kpj�I��^9:(�[��`pin���{֑�*�nIC�5	n��1m��O��U���B���i�Z���ք(���Ֆ8��Q�ַ�!M��jV5�0�ײ}뇧iuŠ$+Նb��=��g�P�v9�'s���^��{�W�{�
�#�#�:Y��-]X������Es��u�e����I��(/�86��D��$�cRo��a�B�a�����D��7��1bի�aꏧ;�O�dSPU����6��6�������u�j���j����8W17���}���և�:n�R�fTG�d
�t�w��d�åֳ���ܱ
eڭ�.���r^�7���}ϊ�vb�!O|g�'�hJmլ�0M��:��,�}��QB�_�'m;�[�<8y�{=9�L��_�<�^4�Z�u�2�K1^Ȭ|�e"n^1�ΠOA?�Ro����n�WnFL�]>�bU�1�Ǻu͋��U/KRh��u+���(��l:����o̘�_9�����˛H�O�6��3K�0�M�tOi��n�PzJ�XhޜҀ�[���g�۫��=5u����c'�2}�:���f�x�;�7#\���}�j����zV6��n��y7�|��ʽIί���j��I��3b��U��z�:I�&�jO,!S�p�Q���n��ξ}h�=�>:3�,]�,IRYRA��<�usч�wC6�
#�
����
�W�����vi�����I#�Y��w�_�g����G�U�.�ޘF3{Z�^����Hߨ' Sw'm���Ч:�z9v0��>��ѥ�$��
=K�X7B[G��g�+6팷�����fw����L[>��2?��l9�B�^�����_?�i���������O������4M���'h���ץ���ژ�����8�������o?����E.�sџ��\��?��u�qj�����yY���=���_�����ϫ�W?�~^���y�����ϫ�W?�~^���y����ݫ�g���#��!����2Ō"��XrBvL�R��������z7�a�M{�C'9;?qg����y���V@�$t��<Ӿ��W�����Ϣ��j�Vz�>	i��y�鸖Ք���_1?��'k"���xc�۫�c.���qC��"��lj\��foN��>�ܯ���g��?_����^:�"�p�+k��=^c|�]�}�(�-��/[[(�gԢE��|��MȀ>WϿ���ԓ��Z��{�T�U���_"o�@�<j�7*���3��";������+�]f�p'�����7��0Ȭ}Gv�/��>j�Ӹ��N�����h2A5�f(��Ɔ*M��싽��F��^\9{d���ǎ<�S��G��h�ʌ��G{��e��d���9�,t�E�恻D�ŉ�4�B��%H!��hK��/�A�5�ۑ���ص!<�Բ#uO]����tt�h�ڷ��O��/+�h�Z�D"�q�4�� (��X���4v
����.D���i6�:�3{����?�����������@�_S���^���x� �B�m!@�e��xt���:k�����{7g�)A~�ٳ���7	<z��q:�?O��n\�eǎ�+����{(T��ީ/|�x���6t/,W���2�-�.��?����C��,��b��]��---r�hn�����蹑�hw<�5� �NЦ��v�W���!���f�NP��~@Ӝ�@�d�-������4Fkg�Ǐ�w�	ٗ�欣C��y1���#B�_w�h���O-�s�����3���3��P<ǃ���SU�B��h^o�ױ����B�\0�+�x"z�2��˗�hz� �Wn�&!�ko�st�T�ϓ+6���_��иi�6@K4WJ������N�����ʀ��˖����K �6����u���
��˗v��n}�L.����V-��B���4c7$׳�	�S�$Mss���_h~�w9�(X~�J�
�wo_�^:���v5��׉9����~��I炔���0p��#ݣl@2n±\���]�9j�r� `��΁^����v�D^^^�8}m7�pH��(mY���e��������I�srr*�oC���=+z�`^��h>���N��ksw�<�<��0z1���9���o{Fgc��F��^������2wss�s����G�Nt�,���{�N��Jhؕ*��!�����֓�k���SGg�ę$��tws��=�+.*�z�Ҟ���ny��E�wWrfff�i(o�eO��g��~w�ݺkԇQ�P�&�?0��p��.�l����w���Ԏ� 剿����u�S .�=V�W\H@����야]����(�u��^8��f���w�%��C�'
�m܀ҾVt7�n;���f0�����py�n_��+ X��A���ce:���s0 ���O�7Q��-�O?�ض�7�<6,چ��L�]t�h���	qC�nn>C�}u�ޫ%|���Z*���ސ��ׇ���S�Q���>3�AF;(�A1Vc5��(����3�m.[�YG��J���=���0E�|�� ���n^|K�r]{A��Ƌ/��������-,��*�$���YK%�8ǲ��hS t,��R�Z�:x�eb�@N�x�h��1�P`���;2zg������_�j5{��U1#��G	ͼ셯@q�|E[���ŵ�.D��9�'i@Z\BV	ьf�_���.���HÞҥ�4|�G���3@y񽯢o�8���պk�:/r�1��k�c�Pn���4-������ U�\����\'�K���{:b�I2W�I�p����ݹ��
t�Z��"�!���.�:u�!�k��s{�S�\�L�q�7`�GN'��v� �����׼nFiM�%�u$d�Tb��;��{��� U3V\B��AB}�?%�
�;z����Tj0d�K��d�U�l9S�L�X*+��z�4����{*�K�
�!���ج���t�-^<��=4>;��0�R�6>�� `�Zϵ����Зhܕ��\k	L���s�S�bF�QpppG�c��^�����f�+g�K����xUcOU��q͢6�t�����斁�
� ��+GUx������s���+�!I5;{�) ��W���F+>?���)��b�E�����.�Ɏ�G3:j�_��ɪ*�h е��Ȫ�D> y�w#/������z�6�ubIXԣ=3���bdx1ۅ@��Q�x9$iה!�مSuuzR���}�h����P�J8~�� X�!^�K���~�����):LG�|�W�/�IY\8����@�[���忴U�?ީ@�{cq�ͨ��*���)�^�yv��[����0ὠT��wC��@����D�!r��M�Rs;�%"�7�#��:XZ�CszΞ�� ����>2���H롍4m��y�� ���(U^�@����{�W� f�������Rjg�q�ǽ�����&��&�L~����+x�T:!�ڹ���(���O���|�Dc���2ю����:r�Hi��f	9�+h�\��s�`�{ (��� K:�h��h=��]QW��?FFcfgeݦB�w�4��C<�s��o��?(߀�N�נ���u4u}���V۪��VPQ�PG�BZQ	(���� dD�Rdoٴ�+��(�� ��^��B
2�)�Y"���G��O�ͽ��9�s�}�����Ԏ�:s|'�u |0�+/��P�@���b�t
�!a�O֞H��+y���kB��*�H���y��CCC��}
��h�#��NC5'	?t'b�<q��Tx���UM���K����!��5�J�QBg��2b���߉l���4�	��K����d��=i�B�脄�{wQ����U^)�6��:?�~P^�~��KM�18a1l<-c��s��B�֢M��`�O08�4k4%����'{�҃��<�&Ҁ��$�G�E����Bm��0M�byP�}�s���چ��5����/�Y���$�j��A-�c�87>�yP��ƉT0�W�b��ZJv�K�zB8ʽE-�̂�$����j	0}8yqee��<�S^�ްu��ya�k�v�� ��t��,��~9���љ����|�;Z�=7�{%�\��lI:�cVou�K�r�NP�z�:}!�8@lM�P�ߏ~�����TȓC�sK���(~�ܢ���zU�6C(������8ޫH�*�(=���hɿ�h9<\gH���&������S|lG"��_����z�,�׏/�{�f�`�Do�G��3��sIr8gOI�����LR?�C�XqvZZZ���|XY��a&��1�_㿑��c�G|v�0����̷^��! ��b�6P�LD��p{q��p�j���p���]v66��(�7��E�A������JRD]�>j*`��Z|Y���ZA�����:�e� ,[q��l����˗/�f*�H�������]{���D�۷og*��C-��Dݘ�
4��,����շbB�������1~JT!G�4��Ign�~(UsI*\�Z��>��sn���z�~p'��O�)mo��:b�w�Yd9K�A�uY�
������i�/c�/��P�z�s$�r���k�Vj%+yi�qC=A�V� ӕ	�˩��_K�mS<�n����	]L��_���r����Y�w=��s�^Z�'.���(ԣ�l��q$"�Z�ɞ��s]tՋ؊Y��,XK,��~��]������8P�&��g�*\�{�KjU�˚�E>4� ����/ 
��٭?�eu��h���/�����_9A�b>-|�;�zӥ��Q�b�)m���]��k��L�ݺu+��n�}�&�t�9�j楫O�2P�|~��
ग़��{�z��(��fR@���Ʊ6 7���Q�s�����v,�b���ήH��Gm�Rh�gP3�%�Ɨ@ܿ��Xp��^*fE��)�g�b�Og,BQ*c�V�a]V�}�ZT��
௮|���{aQ�H�7
s�Q�=�kOӏ���Nī�B�$2�e$O�"�#�J$�5�ķ.�SKR�J]�IQ�:�+m���ŽHZg��^��sS�ǗJ�>���*�F����Y�? ����)S�:����&E�����Vdu�-��u��`��8��7��DD݉��EB�,
Th`�~JK����#&�k���C�c��IE�Y^�S�n�Yȿ��1���"�B��ɉ�٭���R�{\�PW׮�@m��h�B��2������g<@6t����p>QVշ�k�{Rs�1;!ٲ힕Up�cL�����>�X_�#����m=�O��,�L��y?�qh�D ����x�Ȣ���J4^7���$2�3��y�� ��.Sf�s�*�^Ut��T�|	�$� Ԓ�H��Pd�U��k{{@�Yi6 �%��]q�Q�c���R��ϝ(#e撰������	���������ڴ���1z�r���=U��dH���ێ�>�	s�@���!��-���3+Zِ$�a��bQ���i�ROR50�]]],}���ϻ����ފ[��W%:��M��u�]��f@�~]V��m��#��;��y���J���i���mE�#65}�WQZ���!�F�JD52p�������*}���M�H��h6 f�u�rnh�K��Q�T���Ce��R��/gK� ����Ku���s��}��(�Q�˵�"O�t�O(o�&��;��E�] /;��ٝ�%A]�V(Z���ǇN���é��l$0|,��pL��GD��Jzv�FE]����YV��i5^UUe�N&��-o,^�߮��������?���O?��s��ӻ��o�0������[��m�O�*RRd�I����t��x��1�o'>�sݟ���[��ݚ'����V�8��������g�V�6`��n����-��;o��pa�2P������Vp�|��%T]��'���28��n׮�ݐN�U_��b�Ӹr��v1�o��|�-�k��Я�>T>��tP���� p�}�.*&�&�g�1��{�Z͖��v���e�}Z��-�P�إxz�z��<��;]b^�$'�^����l�AN��a\yx����߃�2;��{���A�Y�/.�2����cc��t�R˨��\�6��]�+�cnn��ś�`8T�l�|]wA(oԧM�6�����Y>���	P�(��#9��rVH.�5�a)+�u_������J�]-��]��Nŉ-�
��{��?�)ͦ����	W ���rC�E�Ы�x8�η���{��c�������m�]�֝���K�}�_\Т��{w�X���]@ለ�X'Eka��JVJ��#n����M݆��ޜ�*_􏀳#\�=�����7��,g���(����%�ٶv!�qOd��H��R5f�ϙ��Ǆu�0�z�)~T_@a�b�/�o����Y-3P,�u0g�΃ؔ�o��U���p�]�*ځ+�^��W�돤%'w�Zu�*��9�ϖ�%�m�=Au�y?ڐt������'W��Y��y��mQ�0�It\`GxǪCԄ5i��K�� ��G^��.�o"�n�Q�?9[UU;RkLYj��/�sK#[DmՂϖ���3s�;Kq�o���E�R��=��^�b[ب`�DTq����ڪjk�<��FUr�!\��#
dܳ�m� ����;���?O�6-4�����Sf�]�����T�s�Vm��^m���߼�߄4�`�B�q���w'���V���9P��!� �`>��M

;�(2x��`�b�'�Q+��>�АPᩖUɕ7��Hg�����F�����dCh�]K$�~H��c#�K�w4ݥF��7����'q�+��ii!����.P��}���;-xi���>}�t�i�x��8u�t��ԙE+Y�Z��EK�A�{��Q�gA����0{J�;���e��j�(h1�&�P��}�^�LcC�.�����	��G�v�F�Z�V;�Z�.�*��ҷ��-��Q�]�ioP���E^�cLvgSq�F��H�@���?��3��Ө���6��c�t���T�G�G��s�[�&�G8�zb	Lܠj�8��ꔀ��#%ȸ�6���º�11y����QN(x��ݼ�,P���2�5�b^�!��QG���\Ȳۉs�8+�y��O��m�7;oN���N>څ�?l��d^lb��\�GΉ�6�fbj:�B0^�t���Zr�)��z��X!Wp�nÕ+V��w�T�p	WUF����_�h�pP�㓑g������H~N]'�xT__�R�Ȼ����c�������Zń�ꪠ�"��8���`͖��k.��.�S�U���4�����75�<XJ0��ڂ��U���M��Q����u�{��$��$��q���*`hv]!@�&��'�}J�I6����!R�=��t��>>}+�=5D��6.�јӧO��u*T?�l��+����G��dge�>����T_�2�,H��ī�;��=��X�8@��@��n7h�M�f�vJTQhɯ�(����(5�)�N�x�g�N���]��8Mfˡ"z�k�|�pa6�G���ݶ5Q۬VZ��7)S#��ͳ��%�!�9���~��r���^�?�ª�F%�,Q��� ����HZ{���]�*�l�`�-��J4�f��y��0�j�L��˓D�hY��/�A��M����2��I�|߆Ϙ�B0�@�@eʡ�*�`32�T�uÖ_��9�#z@V��+��c��f�N*��fk�h�7rE^�yiMY���%{����vd׭����.�����/���5��>��!����27���ťK�"���è��S��ۘ=GP4���������WH��R�{2L����]��՘�gP�́c�ȕ��e�
�Tg�֨��7t63�(��{�����"by�W�7Ko1=L�hBcE8�B���WdT��6��f���Bmbх @	���|<۰�ɢ�`}��d yGҍ�+di�/��x������66A~��BL"�C9Q]�Eݾ���[�k�/Š�0�X�^�'�S5[��W06 �4�h�i�M�/��4�E
�F0W۲X"�j��"0+����q\�Q��"5��N�s�&��s��7�̝��r!��J6�6����:f9�.�T(�+�]�G�Q$�<0�kkk7e�]ܑ)w���I���eCǉ����S�t��%VU��վ[�]�o;��~MM�ac�@h���O�~?�$Q�*3Y��� T��/�If�ަ��Sk��& ?Nx[
UF�kJ1�t[Y�b4�ڏlɴ�����ɗ*��_II�g��k�Y�98.�`T���y�d�.Z�W��]!�y1=��{�<Nx�����eBN7 �|p���9/fϞmp�+d':�o�ْyQg�, d#L_ɼ�-�ȶ�F�_����WZ�b���M��w��6|��!��s�ہJ�Q7g ��Ǆ�����'OYʭ�L�	�Q�<a"�-I ��)[b������}�)zO�$���-�h�T�_�N{n(n*ޅq���@���Ċ�s	���"�;1�Gۚ&�p�Q{ ��:놀��LAM�~8 ���+���mJ��D>�\!_�?2\�Y�,�����:�0ݐ�q��1k�GƒH�����A�~�/���g�Y^����m1	U��T|1��r�d�y1{��h[�Y�P���ʷb���Ԣ&~�%���"��)�v�u%m�B�kC��ac3�S�e�3�g����t5�,'�r�$e����[�x�����4)�S���ԏ��dԈL�kz���HB�9fT�)[�lY}���=ᠼb9���k<u[{^^Z�62�5��ko��Ŭxf;�q�3���1F����TJ� =V�-�<�%M'���׽�=}\�_�H�n��������M9��g,JA��=I�⢒c�9ׯ��"�}N+��k�(s���E�ˆ.u���>����:n�q��ER�gk�+�'�@����8�c����Y�ui�� @������NTTT���VJ-p!��{�B7c��*�OeK�D8�o�fއH�P»>i��U$��N]$2��)�ϴwδ6\�@��/S�9���XY�����n��@!�ϻw?3�2����]뷳	g��%'��t�	�l���e�F�����6��b�����������:v�P���*$���455.p�YAH��YJ܋v�O/�^F��  *�D��W$&o�Ci�>W������G��� g��+�b�g�sR�q�+�;��d?rK8�#̑�6>�s��Դ?  ����)
͒z���
B���
���ԥ��b�$�}�����8����:�rEe����+o�@K��w�<e�1��w��F�H�[K]'���iklū�A�w�?�3��J�4�n��8�ɖ����V��mx�`�/uo�뱿<n`f{{{y����S��366�$�,c>%d����<�y�o:�I��̺N�e�چEdV���|u1K�{�33(�5\c^�%���S�\�[�;�nζ݆���U��b�^�� e*���V|vw����l1g}���E���v�eD�/(�f<�t����,��(�����g�����4�HkM(=�>Ė�^`���MU�dE)M�M�d'�)�Dlʮs�Ri?�*�o�<e��O��xrMnG��n���A���ӡ��ָ�M*`]w����u<o,�?e2#(H�ڿ��G�w"v%U>���ƶ�:O��5��΃�$Pt�1���q���$<lg2=ȆnRe������G+�C�
�%�d�B������6�`w��6+�$�5@�,!%�	��|�����dTw����<�L�P�������K���ҒK� �>�P%C�P�N���x���
K��7� 99��M�T�"�@�d�㤚�������,�ʎD�.u�UP��pߒ�zѬ2�ۙ��^�oN�3�r 磷nݚ��t�.��ؘ=vGTq|,d�<�_u�;cd[?�� YJ���7N����з�o�N��dk�ק��8l(9�S�Ʉb���n�0v%''����X�W��ُSy �Ѿ�ϋTZ��܇���q���6��u�,-����D��A�tU�o~�K���1a(\L:���*��n��Q��Aʫ:�3�����ġ���M��=�_+��B
�C6��X��V��J}��X�D�1����m�.��hZ&B�T��O����STY�d���G(o�� Ld}@{��n/�g��Qv����[˄]x'�{=�������Z��å��/����^�UdJҸ�����J���M�LQ����؍��ח������ �l(/�q|=�F0J���Nu�޽��j�$ֳLj%D�M��Q���c]{��h|/�'���Y�`!�����)�<����.��+1�ʰ�,�sf�@@a���g+r�Y��p����;�2�0����ƊɨĆ���	h`����D7r����B]}V5F��܂���x��̻p3j3����=
���Ҋ�)��S�>_���x�� ������7S�.]:@rA�*��^����ƴ���Tuuu�Ν;s����)Uk��l�A����0̀(5}h84���^��bɻj�d��u���DEiʧF��"��#�u�B�p0����,��p�c)p9��N~�zuvH��U^�iܭ�_��2(��<y�V��*u��{s.[�N�k����۷�$>/Po��m��
nE��G
��ћ�R5<�!��yͿN��1߼�;�sY��z$�o{F9X�up��J��^P����[,q�9�Q/}C��F$��U�.ģ"(�V�)oޣ����: ��ǅ�$��Bܷ煬���Z
3��U4�®\��x�&�]�jYG$|}��R�d<� CO�z�+�KP�BTyUT1͌�*��}�63�N�t�[(耱��s^I'5�=Æ��E���;�G�U!r���}�Cy| 	�Rj뷷Aq��o+jKp7�n����#G�MO��W�rr���yw>��g7��!G]��.hJkŶ_��e"NTu�KV302v��K7�8L`�M�r#���}�U�����Dj��[���p}��n�%[���Ե����tf�嘨� �u�T�d��T�
:���Kz�ަ�%)@=IH�e֥��m�+$����C��� fF&�\U��]���D��������^�wQ8MNWҏ
�����
�#�j����US�a�5����5�+���7�"Bh��>,!�@Ԥ �x�=��F����Y-|l�I����l�|^y�eQI"-�п_�Zm굛찗z,�A}}���ׯ�y!�ø�/�)yi��"�Z��ϰOJN�������R�,Wp�nWM�B+�'�`�߻E�i�/_�����7S�}���������?���L䋠l.��xN�P���&L�*�i�kթ�jX>�� ��?��|����q�0sQ���)��="[�[&?v12�]>{���6e㮹�ڰ�-ܰ,N����]��5���{{��΁��(�3�ȑN!{�����n�oaT!����Rp�l��ۦ��wf5�S!�NK�-��Z�|����m�ի��ғ���k��Ny��p������h��
^��l��Ч��8����*O�����-����:o<�L������W����v9ٔ��qz]�[��k?�	��+���P�� an(F�|�M��ꗓ����@L��Bסg5�Џ�Q����U��q��CNQgΘ6AY�h�Jw}no�f�|��#P����h�Mr��9���---�X-5|�K�����,0�Q�IgC&�}CI:��^O�����������x`�*��w,����kQ���+����o���;R��tr�=�$0}�
8�?��4���"�PKWB�{�T��$���� ���t�Jcb�V�C7����Z��ͨ�ZNkO8�	�ޘb�_�)ڽ�Ly�Q
vQ{��բ�&���C�4�[��ǅߣ��zq]����(8�Tqϕo�0Νp�t��������7�%Ӭ�|��:���IϦ����z�yP��yGv]�ɻQ��V�,�5������z���~���_�����}��m��H�%����:C8��z/_8\��t
(l<��)͡pR�RB�Ƽb�k^���6a;�g"�1�SL�]���X��L{��~�e%L6�T�o�E!_�G�I6���@�.P!oF��%<���i�7�CX�A���e����=T����
�j1�Ğ��W���������_p��Ř�;44T>�ب$�.�z�C���N����N�t���%ʽ��XQ��F�/ch���F���bz�U��yp���#����?����m�Z�Z^#V8߽Y]Scx��a[(^�ٓ��u���M*�tom+++5�F��S�5��o�S�^A�bh4�[��}�a����I߯k�>������Ǐ�ƻ�&d[��m9������%�	����d7�&'�Ȝ��E5O\�K�?c�w�xDl�'����o��k��%����.��9];>=��z�jӓ�x;|<���>n��Q���w�6;�KᗟL_�D���������Տ?���b����MI�V��}��g�4prCo���~zqq\y�]�>^�q�~���P&u��yς��֮'W��Hk=�S�c��Q�hr"/-ʂߠ�v��`(�5=%5:�{o���?d�ip����+:��а]�
=��]M9۹�d�(�� ^6��׮]�~:��o;���1&�b^!��W�A�Z6��kM2\�G�5[ʄ�{�V���5u�c�i�'�ne5��'^�� ��"�8Ա\p	uwC��V���Nߑo�=��b�X������	�B�&������q{ł��:j���*�3U-���7�ݖҗ�lM�[�r��8jkR����$.y����)�-�5 ��E͠.>07��dw5O|��%�Kq^!cP�<ǒ@����h�J��������*b���\�꾑�;HS���K��0��K6F��Bq� ��{��������P5>�r�A�]U2���?bl�.�b������%�J2H��=8&�Fo�����#��o~q����PwZ$�����v�q�B��o��+2��{,�IULy'˵a��)-w?!ݗ�&(��b]g�r�h���COf7��u�B9whSr�K��&
�āG�|��s8���'$�W�M���6�� ~^1�Q<f]i�w�P\x=V���#Vb�W��wdKf-���vttXI4��젶���U?4�<�p���B�Ԡ5�2UHiQX,��U^;eHw?)
)I���ZDf�]�6]�L�3=amL"X��n��Sb�L�W(�f6ct�R[V?	��	�:ګъl*J�toNx�F���]��鳐�b~���"�C���1:��הK��-^Ê��9�lb�.`63 ޙh�fwZ>����Q��2����|�&r ���fw]z���PC7��e��%�*�aR�����K0��PR�l������c��S�4��+$t�i��{�����ii�XܻE���\�;��V:��w��8ө&-�e3{Ɖ>�E���&𡜥���P�JĽO�=�q�˵�'U&G9���lw���óٮX۫���ϗ��
F��1�!�h˃H�Ȓ��\ID\	��/c�V�^�L�6[.є	V�!>anT[`����
[�*�sTvi��^د8��Q��q�#��g�T�=<���ᙟ�J��i�s�=��.fff���`B�Q��h�	��-̞��l�᫾�Ř�Ը̀	O!Z.QѢbg��Rg�,N�K��eq	��ϱ��U��~������v.��=���B��#�"E�̳����z�~'��$�1���K��JDi��W_�Ut��!KXխ���s���N_U��t�ҹ�ր�Y6��w�
.���mO��ɸ�!��kI�R�M{��P#�G
�H?�	��~�#a�&�W[�,lk�]3�Z��8�Dcj���BDQ�� MA��g�G�!��r��!u.ٝN1�ɥ�EQ�H�ݻ�������e5ڣ����g�N.�5�(����\�5���Ib34Jڵ���Sؕ�5}�P���م�d����Q'/h�s.+/O�ыS}!��R��j�����Mv;���m>q苢�y�a�ڏR�;����*�P��Z�w@*H�e��`�u���� ��Ѱ�7R���z�I��t��o$�.��r��C����v����Q��l��x���cǎ%��IJ`��1�CqS�u|��9uLv43?�w���x|��wX��D8���E���ܾm۶�h� 2�4D��S"��)�"�K����6�����x>)z�U��ʽt�1k�DԞ��ڳ�7}��sa䅸)ϯ�1�AP@=�
���Ak^=����Zo{*��G�leU�t8OQ�p����:��	���zf��N\�:��;���������ٓ^�A����r0T�n��T��C�^�0��Spir���%{5[\[�7<� o0�
ތ�5���R�־K��e��k��f����ɩ����+L�+Z����|����aެXc_���Ǵ�v�{�(�?���&'���kW���V�_��[���*���)��H�G�J�=/���	J���F�9,�1�[�nL��k�-�my!���ՖS;��	5~J�<ByP��L(̦8S�#�0���-����b��5����K�M�������Rw��5��Nÿŉ";���8h�3��*�+��fW꤀r��IPU\�r�{R��Rp-���ݚ�+��6*��<�%��7}�D*��G����X�0�KV�Ă ;�hCV܁�+��!,p�UU>�%op�^}u�� E�@z7a�Ժ��{\y$���>�ە����C�#G�*SRR"�Ʌ����n!�篢?���KC�_�]��ܨd�sNԻ��$:����+{�t%�{ʢN�3u�Ļ|���*N��\y�֘������K�y�fS;����`�~�w��З�x�ak���l	)|�=(�}x��yL�M��Y�I5
=���{孧�sv�ᆊQ� �����(>�����(�_�jD�!���52��S�u|/=�U��v�}�Z;������\�:ȥcg�V��� �Δ�%_�\������� �i���Ww�ګ3�5��ț��	Р2�����{����:YT�(�_���J	o"2��íڑ]l)
W�za{� :�PHΠ���s�5/���5���0���đ˩�cf�:��&�٭��U,*G*> �r}���P��CV̠QP0o����T�r'7��2�N!c�N(��._^�P�B�{���T�����L+/cם�Y�L��������Q�;G���F�9�"���L}����u��?M��^�	p�����M���G�G�$xpE�4ژ��0p��o���M����,wq��
�����ׯ_�K/~����\��
�U�&��&�cؒ�5���G���YM*u�}�U_*��K�����,D�#����4�ݱT�>��e�O�am�3�E�6ox襔;a�os"7�;�7�%�;���i���?`K�l(�c����z�t-�!��a���	ԌQ��m}�@�����A[j���E�l�����a������d���w4��h�_-�F/��]0[RC�U>E�{�߉���wL	/j��rK�޳�|r�Co���"�=o{�j�ʙ.��+��(\��݁6��.��%�R5G�($��;4��=_nrr#�f1���c��ΧJ:]L��cTMA^�p�p���9K�=.����S��4�J�l�]�v����+��wSݸ����Z��r_�9��<\���ˬ:EvH،57/Ѻ ۬�~��	�"%�-]�rd;Ⳕ^t�m8�4��9���G�}ZK���N��ZY�=%ō�9l�g�����>��J��S�4E���Sܔ1��|l��=>����0�*>?`иL�FH���t����c��*Z����P�Ol�̥���K��չ����n��V\y�&������̣��]oo����K�0kr��?<e>��YxM���dx+�CX�$�`TԻ��Jrp=�� U���n�P�X�x�l�0��\`b��U�D�#���ό�A.�ߌe0\X�Zy1ќ)��0��Q$L���w�$����OY��y�T��+ߎ��L.�hgʹ1_ߵ�[O�U	{��I��2y�}¢��v5["W���
��"���_��aDp彚-K�x�m�S�x���J%ͮ@�����%�r�u�6�^�K�u���!w���dC�P~U�����Iz�H��<f�qa�l3���\�Rzѹ���}�����-5[V���g�I�<Z�����؄���y��L��B�HW9�F��ֈ�6�*+f�;eq��oUEE�L⚟ӳm���z9Ӄ��D�����5�~z��5΍�u��)U[�R��
�C|L/����{<���PK>ڈ��m����֣n�Ѻ �\\k�������X=���CU߷#����@�@F��#�4Bx�az9p0���,_����������)�E�e�R��!C�!t��Ԡb��v�7�i�@F��"22�JN��v��/
�_(�����w9ò�/����ɬ������Ya�W�i��K�Z<��5a.SJGf�w^%�3a�;v	����`P�.cK��q_���%�8�ig�+�u�R�+�(26Y�%N��O�c�>��lieG����$F%K�v�԰߹s'�(8Z�NLW��)�g�� ���Y� �W~u��*��w{ ���PP����Ӈ����3>���r�l�UX���f����/����|M��Wrr�v�x��w'-����q���?ƒ���b��C�?7�t�W�B?��Ç��>���X	�3��wym�{�ҟG�܋��r.P� 2��〢'��'zBQ^�[Cq��,V�����^,�3�cH��Y�~_�z	���#�H!��&�H�Z�|l3:}�����U��Qq�>�+R�%0��V�x�O�(�~��*i@,���zy��"���%�X8�������h��\ya�]`�y%�k�lP�-�͑��:���i1��\g@�|C[�ʣNߦ�2eǄ�Dz�F�]vv�7�K/�p������a�"lQ�,�c�l�_�}�ї߀ĉ���Q(���j��]��xs�7?�5�
��]8��)}-�кn��Z���q��T�H� ��vL5���T��ܣ%s�OԽ�،W�O�˹\�ސ\�~O����9���y���o��F�p�pG�<�'��~l�y�EQ|S,<�}LOV��>|�+�E�F|�/�އs}69 ��C(܍��.
�����O �he5��nJ�̵	C�D)ަ�I�/`f�t?��w�M3q���Fe�kh0G�'�/�{�:�xM�W�o�K���H���,ta�?>H��&�|beU���8�u��g�S�
�s2������*�	T�G�-��D�)�X�x���|�Vԃ��+J������I���$X��;�
P�W+M��~�0ѹ��%�i<��u�]��e�'v͜�ξ����6���hk���~ژ=�`є�W�4t�@����������Ŭq7���C+V� E����q]�S�vO��W��IT���(���`�M���a¿���1���Ht��>R\�B�&�jP%R�b#^=��m��)Ӷ��qG�裱����Y��j�j��%�;K��k.��
���+�%d�d2��U-�@���	��f��,���j�����c��}Fs�q���>3���1����9�1M�V�+[Ҵ����*��
��Ԡ��7�^�!p�XX�&ܣ��Ɇ�{HE�}�kX5~Ёf�R&�sX��Q$��U�UP�� ]N��1��''����r���]��j��jN��
�����\v
�~�����n�
��(}��p#�P9rs��zcQ�>�JgL����E� ^����ü����� ����}�~D����v�l�|�Ԯ�v�'���N�;�Bx��ǫ2�����4��ܦ��T��&��dac9�}m�K�{�F+�`w�g�"L��w-z9DD��� ��ki��þ`�#m0I`�I��|�q���*G��LKk� �;=�fl��ڞ�Y��E�/h?�q��$9��S��K����hqW�v���l�/�|2�ri��6~�$����5��IK�*K�e\�������璓#�J�ٜ��̘r�#N������G�?�m��w�C̙���8�-����#!�:�ad܃���ӧ���;�Q�K�洽mʿGl�.��y�-�!8e�Q�� �p�fZ�O��}����0�z�^��P�Dq�
���/4wM>���0*hK�������.�����.mN�� ��hm���ҟ��k�K�GA�?(��l<�-�pʴLRE�r���MÄP?i*&�q���E,�MҞ�������5�9HP��P<G�Æ�(D�Sl�wSff�1,N�VO�w='g���� ^^|'�V֞x��y�C���9�VU5y}��';�X���a�J��C7<#/��P]�����H_�������f3Vs`���bʡ�h��ct�����:�+O①������dD濫L���0����|���ޭ�?����h��}| 3^�,2�M�:0f��-͕JHuK�A��k�z~ۇ��=�l��_�x�lԘ؃
;�>q���$$+t�YZY5�1ˏN `�����!�愨"$���[-F�VNڪB��S6�2�g��Jh.~��E�lk����{���i�ţoG�n&��~���n�;*l�\�9�M�bH�ю���U�����B�~z����=�NE�ǰ�/���jO�����?#NY�.]��ܘm�Հ�y��!�NX��8��$�1h~o��m��	߮�;�����u���X�����/�?^�v��L���e�Vf�H-]V��.���3su�Vtj�����2���{~������?~{�����_|�KzV��V�>s�m�ee>	^v���c��n.��ߏ��T=�v�knk�P�(��� ~��^��fS��Uq立�w|��ӑ]���ں���͏�]>খD䄗mC|�28��a��CZ�������/�������U�Y�Ϫ,�֞(��fVk;�|j�mc!і����^)(�i*�9����t=�Ws��!Gio��LII�(��d_�������rp��Gh�ϙ>�~�d4���zUdQ�����נ���]wtOjߟ�������0�TƥDGK��e�e0(/U�v�c�F\IttMϴc2�@]əE�.uq���F{�V���[g0���k9�@�M���{B�쬛~��L�řk]������F7�ÄB5�#�i�E���g�J�n?6S]�Mx�
C�E�Л���י=���f�X�D&*Й���Ꚛ��U�o�b��0yu�ʲ�\��UTT�f��t�f�����<{����1�m�D����0p���=N����@j��n �m����7�Um],�����w�.u�Q+�tX6o9nta"�d��rI�Z4�����\���,����2"}|���2=B������q���awV�=>�	n����r���˓��O@�-��gV*�:�������c%�o߾O�@W��MN1/��R݄�M�ԉ���������1����ze �g�����N���R ����0�"���<b:���������w_������cD�g�����}���$h��ߙv�/%>ř�%�%0h͂�a9F[f��Q+���5(�rZZZ��X�ƒP����C�
ʥ���wy�:��/e�,3��Fe���~��̣å��C7�S��V�Z~�d��vZ[x��(uM"Z�j������ $��9E�8W��qa�8�j�K]�݈}����������#��,�R�i��Fmt�HϨ7r;*@��4��-�k�]�,�Μ�7*�s�2u�S���r�ϛ����|��k/bE���s{U��+@���02$۶o�o�0{����L�2�=�ퟔg���X�u;��1��s����H�AT@a#@%���n���}��w��\V�M7��tC��2qɖa��ŉ����wE�2VH��i�'���ݘ��Բ��V�dե�,j��ӎ
��eb��ᗕZq�z�O 
L��0/�n�����'խ�hZ}�D��5��Q(�dPn�|i�TR�Ǌ؇����/���з�?��{�`�S�� :wxl�֓����87�D��T�_"����f�};�x�\�F)�hխcN�QeZ�ʼ��� U+����4�8T.C����;`��&������:t�`���!��[i����8O�R	>L�4���ΝC?���
�q�$��Nh $q2��tl<�ZDC�%��^��Npsr��HVK0n�1_W�_�	��4B��p�f��U�3]�=~��핽w"lg3��=��t�G4�J�`�?�c#��#�Ba7�Aҋ��u����n�r/�����`�6n�Xr	�
����g�W!#�.�.S��:s�<ح� s�3\v�d4{pՔϣ�NNN5��6��M�͏�Q�'������X��p�����S���+vM����3�%��(�^�m"'���*uC[~��y�9����E�dj�q�4�ٍ���r֜�0+�N.�h��兗��g��R2�����x�B�����W�O�N@���6��
Nt�����95��c��-��JF���9ȃ�K���P�y���:�>ʑ&z[P皟��߹��.ch5��R��酯l�v@��˟\g�<!t� o�`�G�.�%oRg�u�ԾlVK#Dw�W�ð������@�˺���K���#����s�D���U31SLe<4�TExE�u�ԫ��Zt�<<z�V���q$�<�R9bQ��@�@���Fm��BZ��n@iAJ��jp�Wto���6���VE�I�,�؈�cޓX�OW=D�����+���$x)���fy�y�b�a�
�;���IU�Cϣ�d�Ӻ8QPȍ1=�y�pa������zGN
�3�a���}~�L�ޘ�8�6)�u�N����R�\�v�֟y'P�e)��!ޟp &c]����� ���Zv@|���z�J����V��,Ѱ�z;([��:�4�7�~�ŉ���#@<v���	D�ƣ����|��Am��cr�A&~�ώg���yV���ͤ�P��d�P�oV(�Qv�7~�	p`�j����~�nH�����#>y�|�	��F�K]�;ɭ���"U&��h+�(������N�&��O�c.x&3��������7�t�BV�Z^���K�*X��'_)M���5��S����\ �b��+�l��&����E��[2�	�D����	��{č����������F|��0�?R9��~�`g���2�����x��) ��2P�h��$���1r�PX�f����?__�u��`��>�Њ�Oޛ�K���ֶ���Yih�9�}�o�хGG4[�P��2��~�/'�\|����Ka�R�������]��UUU��~���3�X�8;�1�^�(f�q���K����ւ��fc�}����t�A%�����p>����i�S�Oz�MR-~�٘ġ;B�h�������P��K4竇n��ރ9[�3>�t�X���vk���. ���� /}��
PoB�D�0�9���^=�e�`��9X�,�;6��mx��v�����%3׼�Z^��� �ܢ�u?|�|?�i��RSS�/�i��Q'e\ڿk�����)�{4!#�]�i_���.��:���a���{?���=�"�#KN� ,K�0�^�'w���P��;�-�[���)�C8����yv����vu�����n9��-�v6O	� 7�M�*O:��*7f�Ƃ��#�z�G��?㧏�p+'$����L�_�9n4 �h<�?��xAg�0�<ί�0g
�����5�r]V�� ī����� b'�L�
u�>��B���G��Ї\t�z�|����y,���UgMf#Ĭ�-�𽑁��t�릂�J�'������YL{��0|��s���9���'+��v�CQ}�Y����|�rPr��\�7��R�k@%Ow`��^h�� ���]��{�M�$�"��&_���'W>T]]���$
#5J������.u�$�vD�|d��
�qƑ�揭'�}gY��2�ָ��Y�;(�|��0��ɬ�*#ѱ�I�b��ə�����K��u��o�M��u{�ۨ+�@��-I@�ː0vFQQH��-zO���Z��0��Щ{S�)4�_��Ϳ�<���i�/����PK   u�X]��  A  /   images/bad899ba-ddb5-43c6-9f63-2d962537fb78.jpg�ygT��� M�"H/

R���.`���t�&҄(� R�H�r �8��H��[�B�������޻�g֬��z��y�={�5�i�p�H�P�� �P0�;��<�yVfv6VvNa.΋9�	^��������RPӻ��|WYJZ��]#S3S�ۖv z&��4���l�l��j�D���?7Jp�<PE#BKs8w���"��&����4�6�5�s�t��癘Y. �hhi�������Q{©} �Ez�+
:��O��q)�M�~^�nu;�����J��#��/����_�.!yCJYEUM]�ֽ��z��F��-,��ml��;����{�|�.�}L쇸���i�_�f��(�YR�WM-�^���wGgWwOo_����5=�^\Z^Y][�����'�98<:>!� �4���x.R񜣣��c�͹�:/��_Q`��3>��tU��y���߫ۙĔ��~�?�|Y\y���?��E�(����o<4�JKC0ڋ 8�����?��f~���� �	L���禸����a�䦇�l]�����z`%>���T�^��_Q���Wcq�FwO	���8��R���ՇY�1k� Nπ�"v�[K�3Y��ɨ-��h'�F�x"Y�4�+�;o�o綀�5|yI�Lk�]^�;��&4qv�@����bq�ip�'F��y��O>y�h����S"���>پmYc�į���(��V>��{�O���|1Lu|�� �Tg�������'���`��N�Ua��k����D��h����˼��{�
Z���!�~FƐG_�����k�<�K���rܠ�*��E��������	�(�w����:%�.����V��Q��Ȳ/2�܋b]G@��;rv�WO�?�>�� �5U�c��_6����{9 ��{��$H����r������l��e������Ѯ<U]�U�M��]%���tɐ��w@�/��N{��b�}��W'Y%����S���8�n��×͡��'����
����	��^*[n�'C�ȗ��ْ�yX��t�{H�I$
`F^3g�Ī5�BB��N?����q/�,q�)@��=��X4� ,���"���}���`��>I>�����A
P�jt �>�����@���d�=�������@���.�4w�Q�:1-h��5H��Mwإ\�_����p�������P�
���.������q�VB$M;�n�{���!�E0o���ٗ1-fKU
�a�D�<KT#a��V�,���^/�(��Ρ�B.a�rt���iP�tt1�X��;�}/ �yT:f�� 9l��8zzj�j��Ɨ̩Ti=,�#�^*�z"<�St�Н܇f��Y��-�?���A��u�v���$�v܂� �
?�}ۿ�;�����NiZf�j@1?�s���.���P�L�����F����֋QC��|U�%ޘ�9����z�I�Z���כ�L^y��J��a���G�?!=28S}ᭋc�כ���#����Q�͙��m���J�o4��J#������ii.t�~ߞ\�~�`�~ �92�|q��NM�c�F*��+S2��Le7�a%��3ϓ����f���$Z{�d�3
p��7�ؠY���z�Ω�}c���.��V�7���.?-~�`�uW|�v�6JRmn�s���vh�/�H
�*`	l�+o�4z���3[�\N�����i���>u��g�%�t�F���M���k�O��|��V]8q9&�� �n�m.������9�Ƥ�>=�\Gx�&�%Sw|z+����EގvX�8��rbsS�Y� �� ��A���8��� �u�b����k�Ц��.{UG���7�-�y6��d����F����ؠ�ǧ�|C'i�񒫈�\����Mwド�٥�YJ��&�ڣ.�c� _�2���7��o+��Hl��&Խ-9���Ho$�p��7gl��)��%��J�E�$)@ 1���r'�h�jo��y���1x}�W��]�����%���˂��L�U"å�(x���u����Y )��8nsr�ǫ�K3|{�[*�Wk����������a����/.�E�+r�,���4�Z��B�~:��{���h寙��������x)�����մ�RQB42U�T�i�K~Rwl��u-z����/��������K��9��?O:��~Pj%O<���jz*��S�lF�F�h{E������m���L��Oվ�Y��L�=�l�,>U2�l����1G?C�hE#��[T�B������5[7��/���K|�R����$P Y����2��gEEF䗾�KJ��'ӌܹ}�^J���S,�����b������o���'25R�6|V��#�7L:�j��k�b߉cOn����#7]c��s(�=cA����4i���l������}�n^o���^~1=f��d%�o�Z>@�	� _��#��n��I#�h����9���C'��(��&��ChV�
��y~9`����)�SQ�\4yˑ\�w����I��Ѯ�)�c�����X�N�N��GmJ�(��yB�����b�S�gǖ�kH��n�d��oIvN���l����w�y�>1�n>,�����ܝ�5lr�b���mX���^1�DF���%�&�j��#S0��P��w�l�JE�h��{1�����݋d���v-?p9�g���� Y�7�����9�͡�#�����p��W�r�}�����η��E�}��I[����k�9�;��o������8uYա��/Zۿ�_�4�����S��,!�hB�/?bO��E/�P]}�k������q�]@�H�t�^�e>��θ�g�!�I풃a^ٯ.���٦����*V5�R �dՓC�γ��ߡ�4y6�<pb��X�4\}�X���~#���w�~��
a����e ���@����r� ����w@`�=W�`��#�Ŀ�t�K��u���{T�4�G1-����:�ܐI��veԸ皑��^H?�\�`�AL`��A�jM��M�T�����ܭſbE*9D*��O��V7�����[;�U*~�9)=K�C�h!�J!#�����8��)_�-�q��������gϕ/!"
a�J.)Жy���+��1���e��)�ը54�q���
)�x��
��b���f�q��%NA�!'&�O,y+�ۺuzjYf$xMe��%�Y��@�%#�E���PǍ*3��㋎J��O�'&�жkhBJ!S�r\�_Ji��ZB��l)A��l���ʘ3������	�~R&�F�?��?ѷ���}���@� ?��>@�XL�Wc�z�����f�����,�3�o�	�x�ƕ���ޯ���:W�3��/�C�]bz#�c�?����� �'I�U�¾X�X�i��5�i�b���U�"�.�08b�®���Y�/#��r63�"!=��U����Dݏ��4t�
o���Z�Ԥ�u�T+�=Y�W���t��R'�Z�7�A<.��멲���]p�c]�,X:�'��������oD�[F����0k˵}�}���<��4��7,bI� ����� 1%>����H`XO�d�J��Bqy>�:�2�0�b&��O��jS q���O)@ed	�5mO�#�܎�r�����c�+��ݸ�O��t�E�=���<�;�Y�O�$�qeg%N@��A�QK��T��|�d��2`�9�Iz<�[_�":�0Y�:��m�(@4��Z,�*F�*��Np�^�q�[a�;1M~�3�_�|g�����]f�w����Կ'��w$Xd:3��x�㿿�g7���S����_~�ۉ�ݠjk�K�eU�D?V�~�F�O��y��^sv�p������oڂ˚�y���sϷ�yy�WC��G�lm�`X�7�:�2d)E���k)<I�S��K�j��]�d#�f�jW �3����7:�9�x;m�>�#��3t��M��� �}xN�P<�7/����jw4s��:���%"��\uv��ͬ�a��'��zQL�Q�T�9��(O8ƳJ,+@�`��r*���q�W?�������ص�R%��H�Dz�Tv<�[��r��L�����^`�y�v*�}'U�/|G��O�PK�.s����J��"e� u�����[�9��1���C8Orl���rnY�m�>�ߺ0c=[>t�T9�Yok$�i@NK����"x
�k���~P�������3�����q2�-��F�������Gm��ڏ=��?˳5�ߤ1G����z{Z|KJ���(��6a�'aN*��,�t��b��ڷj5�O�Y/%�(�(�I��^�d���g�}S�'#���?��ɿ]9ywŉ.i���\F�$f{��Z�{��ր�!�F���De���k�)��B .���J�8R_�hu�_�� {�s&�)&���:�R�/�%%Y�[Yĩ�X���p�~s�ON}�9�.�U)-��[��Pގ	r��'�
��έk��iz��[��wR �	w���?�%>��|S�'��m�>ăƠُ�����xH�j�K�9��I�������ߙ�ǉ�Z���.^l=�d.��eGBρ�7ұf�`��V���;�q����n�iI��>��'U���ct���l�����/`}��t'����Z��O���}	E�����V�� ٿ[*���G�#��)@�Lƍ�ƳE��.7F��GӖ,���;/J����Y&�G��9�@��ی��*�+(�/��� �mm@.ـ2v�Jȼ�@w��]�`��s�qj>��ޡۼ��LA�\69RQ}Kـ�u���j�˱ػ���AV�ݢ��TO�W`�x��.4䯶�Si�G�K�����
ߓ��_c����w���Y�k<Y}�	�6� ��=��́���Y�x�󰱦�`B��l����Jfȸ�=8,%O�c5�8{�����;�F�,_�	����5�5���.x��?+b1�L������)*���Z��"O㤓�������,�Ù�$��h�;��[g/��©y��z�M��JÙk���Z:��5	��=�(-Q`�����^-y�p=��F@"4�!�~PѢ���r���P�6P�I��d�r������8���X� ��E��k|-�����b�������xҐ���b]������B��B� {�9G�\MM�,J���π�"Z�������If:>�#e�Mq	����Wͩ��������k���wp��qv��]>,������7{7n(+�mY���]К��G����a㐲�@�S�A�6B����~�@`]����&k;�؍�ε�B�*g_�8v���rh������ׅƔ�ъ}I\�k������8#bN�Q�[-%:�nh�\�h?�B�mY���� ��x�#
�`;n�/��h�7WL�ڠ������Y���w�w�5�(@��Q�Z�y
0���B�dXG�j�3`�'hi�l�䙭z0:�t�{{L�9]*���#S�~$��)�֮��E�#������z�3n�ьd
:{]L~ç-�zep���c=bi0=FG���
��ij��r���\q�}�Ɠ:�lѮ��&���:�	6�!u���aON���HƯ�Ht���Xq�YRI�9Ţ3ngU.�'�v�'A��>G���?��g��UO+n�v�**`��i��Q�e���2�6��*{��@C肎��6�Ǘ����{H,�xF�?�ƈ&;lDHnim�x���AW�$I��l�K_��*�e�ȚjE@�Y3H("��i8�\M��D�� �{��0�=w��
ӹ7��Z�f3U$q8�S��{I��t��'����zt\9��2A���yu���:Z3��H��Do�,�:Ӥɢ^p5iys�����h�Zj���نGs��N�t�#�Y�B��5h��E�B�y!�Ɏg�_FMx�:�*����
��T#d�Op�y5u;��Ag(@+��'��l�� H*�R�e�z�{�#�YE������t6��{���g���?z�r�&-1��\�n �J�A�!�]�Z���*b����vI��O�T]�q�����-������)�Eʟ��z4�(4�� � a����s����>U�۲a܌���rG��v�ہ�}��,
�?�؆*��/�YU1'!j55�i/QZU­Ȇ���Y@w�X���X��o];��T#�����=:o�~��D���HU�ܮ�.��+u3�ű�M߽�[ԃ�D���O�֕t��Ŧ'0`�J9�&����m��=@>���]��!����ܕ��/�5�ɺA.Ч U?O(�ۊ���r�S�V�� ��`��a���1S��.�嚎.��s�/���v�p�O���>��Al𠾤���0�4A��Ґq^� �P��b�`�� �7�XJ��#�sc}rAx����rf���^,[Q���BO	B�)�_�4� �+~uKų���#������}�_�k���C64*�Kѡo���J�� ���QÆD��
=놋'˹V{��Wk{�ZLu�7�#o?I�5ZR�����3pq�cq�`PJ{u�e*\�SBɔ;EBl<#�
��ߊU!��T�m�MX?���;ǵ\�^���������\�M��e�n�2y��<��~e��h]G6̆���2?x]�0D�(�O)�T�F&����� 	d�43���H�[%�"�m�G'�)�٬�̸�� U��w�˺_�ϻ��[�=*����2,�
H��Hz8�¦+P�$a�HM���:rx�"뵷�՜�G� Ǔ�a}Hִ�[��jR,�^��r�Op1ܓ���/�zBa�ċ.u�e�X�m'�����۲9B����>|#��@�J�.c�7�M���9�=�o|���k�g��]�y��C�L~�3"�q��×�e��C���V�:�T��w�F��iT��F��TWqwy��>�]!a'�;��Fi}��h��.�38N��a�&
@����Z�D$�4�`3����N����v���%�V�U��Y��D�z�k�����J�����S\rwbz�9|M0"�?�Ď��d����2�T�u'��3EF�>�9��V�7uR{����%1Og#�uҡ�s`�=u��%�d	{����-v�Տ� ����
��9���%�&'�1����s}53�~���?g�ϕ�B�#��wϾ
r���ct�������>�����g/��G�")@�ք�H��;g��d�ڱU�7�7W���K��z��S����G�k���x������@��*t�U�,��m'�d��t$t�v�( ��I����ц���霫dn�aI5�V��P]-A��=7���7�PUx[�
��<����S����/�( )9܋"�䬷�&��$�m�e��j��ڊ5Y3nm�)�z[CV�=���:�D<�\N�h�^�T�xXE�
d��8a��_E"@O�rq3�\`�?GQ[��%����W������?��A��ت2[���R	���hAk�D���޵ Kb�ǌDT�6������a(�J�ݷd�����Z�s�m,^�V����_��X�ckh�w*�i\��/��sѴQ#&�SzRR���z�.����?� ��PK   .{�X����<  �  /   images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.png�YeP^�'X��YX�C�$�������;X�ӥCJ�E�nI%�P����o��wg�93�g���͍��Q#1����H4ԕ���v����NI%��g=�M����z��~'C�Nzcw{��K,~'7o[��K~w/���2���4�
	��bz.k��wx;xq������[�����H�S�^��jz,��D���K��
9��+O��,T�"K��B��l�&�|?�u���YTT��1�2������3�a�!t��ư:��4��ޖ�[�\È��9�s(&�k��������]7]�ǃ�A�})$�%y�4�?u^d+�O�����k�Q�b��쫛�'�k0��b?�����ckJ�,�}��+�Kd5��Ҁ`͜�FJ h֊�d�OU�Yz$��D.��Ff�I�g+��\
1��{F�rV�7b��R����	��b~���&()�Rz�(����,��0��K�JQLD�9�R*H2��D��x�щR��㷸6ΞF>��U��a�q�Z�$Y~2�By�'6��ZQ2��`k$�bI�������p{]����1 v��X��f��2��7m�AKQt���L�;�{�Ե��h����czBSiH�D��!Ź��[La�����;˅x~\�%�f��T�ϖt��ߞ��ǩ��o���m��2l�f�:������>bE3^
�{�V��(a�r��^�.�L��)C�5{ǌ��!�?�W���ѝ>cl�4'�p���؊�g3+��G+`t��n����^V�L��4�}�DV����f�Pj ��޲dq�"m��BP^���[7�B7�\����7�:C6�=���\IIvZ�\����]�������
v��vG�,l���=?L
�0R=ƣ�S��8U���
�d� �?��>�[Nƻ�1���sLP@k����<�oD��ZY�U�\Q��q�\h�]� ���jnB�uk�I�ōre���<�ǀՉ(��^��/���3HԞ�b�M�-I��%+o�.���׍"K����hFt����}�a�����iiC�����7}O�6}�`���^st���Ƚ\�aB���TC 5a8Ԉ�,J�s#
������#�H�cS5G�|}�2����6�B9Z�I�&*֖_:��-i`�U=�1L����ӎW�o���p��<D0Va��qC���"X�_�/���7��dB�.���U"ST��u�(�;RQm�<4�E��c]��?Xfa 2��>�זY!����]��\d��d���9!ɐ�*�ѯ��o�9)�b��w�iF?a�
� ?������wY[X�߶:^OL8�-"+k�Fp?�f��M��]���v.Lع�O ����pL��g�,��&�L�릆�Qk#�C�]�g���*�_������N�F�G���i!U.�JlT��r��MDX	��J�L��p%����ƻa��k�>_� @��$��i�G-���_e|!o�Ш.�x�I{�XS�[5V�<0��`�X
�	,��RԝD`��6r"��Ya�[Ǌ&�+�����g��������^k��qBT~GG���Cޫ	�7T.�%=�Q�k�~z���_ǣ�u�*2�z��p(z������L�zkļ�Ŝ�#�����
e.6�$��O����ެ��	ZQ|��"Yz�	Qj�h�S������.�}3�����E�i�-��䲵��0MR;���<]Rd�d>Ɩ�c
�P�w�����ЂD}���{���zΒ��2�R7����;3��������w����9s���1����g���glS�87�*]�y�C�|6�Gg�4Ϊ�i�j?�3��i�9JuxT��f��� w7k)��YLY)�l�#1Y�D��u�-���*��>��!�@C��)�h��#��V"��?��Σ�d�?�r~R�S:��%�{m�F	};��Ě�c�c3z�}7ܽSa}��g5C���f�\Fr5�
�B?���(\v�7�/vI�⧥	3bb�^���������"&��,u���(�~���QD ���PJ�L�^� |䵖>L*� �'��Ԟ�URң�Gїv�Z����C�|2&.���ܮ:ۋ@�UX+�fG��Dn�m;,�oC�ݗ�{��/�p"��I��b��`�Ӯ�[�nXK�7a���!�WIې��j�*����eЦ����V�7��|i�ܴ�����фRO��/ţL��B� M(S���~��GVa>#u�����ӕ:DD��=�r�y� ���zi�D�� �Ò<� �J��it�e��т���+-L�:(�I"bZ8/�{�F`�i����1�j+�+!��qJO�B�ZM��ww/��-5¸��D�Ulv��z�2��!��P��G8��ZT���G��4����x2�#=�k4֍����O���V� ���pбe�ˎb�ǧW\�0s��<���{���Xa���:T�i����_�N5N�(��w�?=fd�w�Ƒ�ֿ]�|8�j�4F\'G߮�xً����a]0j�*�By�����@��1�L�����
?C~r�?���n����j�{�?��5�P�.G(]�8I�i�*2F5{�#��]�����l�X"ȓ�>So�&U��Jg7�^��GMd�`�@hhw�6�;[��1��YZ1)͍y���ǫ�q�l���S��-tMM����Ry�_�hf��Lf2�����4L����I2]�2�c6%�٤լ��s�ha�Iq�y�)%qP������ڿ)x��%�Զ11�x^��Da�t���`���x��H���;��c��20q?hv�4R��|�A��TK��4�"�����[������h|��hyg�߮P �J�ߞ�=,
낊$�\x����k�����W+Ԇ����(]�b@ER�J����������/�X,ү��b�	x���Mp�E��L��q �)TTlٿ�+�RC���a����"�v����.��66��϶b#���X��yNı��U�j4���ԥ�9���{I/S��Ola�A���}��Hԣ��Yg��5��p=8�)w�%�c�B�xyRLu��\5S�I=���BU��wْ�d���>�JC��_[s1�p�ˮ�(�Mkd�*k(x`0y���ϼce��"�JrU�_�6����X<��?"����ۄUD�Y��k� 	|a�A/�zЛ"����&��45p{�wo�7���˗�-�Y�63�n&�\�G)Ekq�#��b��S}i(`�\椨k�o��:/�'xL��.{���ǂ?���(i��p���R�$*�S�e��ͬ<���Е&9����d�*+Z�\���5�6)+��@�O�>���#�a�5(�}��?&���F����t�C4��p��Y�ݽ�0Dwdz۹��)KNؿ�&D����Y.����ʊⱢ���=J/�
��S����U[7���-p�AR��@�r,���t$MS�����XrZO�?(`)�֭R�H�i����]y20�EU"����=�Y�Xܭa�q&i",N�ɵ���j����]���������`YG��3��ڲ��*�ػ�y��~{M��@� ��:j?Ď,�3��7�頤~��1L��"���M��!�|'2�2����ʩT�۞meIR�xH����J�۶�E�Ĥe�Sj|j�݅������ �M�frP������n�U����<�C����]��@3z��Z=8Olֹn(�Z��Z����/i��C� �dݍ�N�>$��4�yp��o�rO^Yۈ�ԻB��Е�ސ�jFɉ��Ö�VYw�K���6����wYg<6���ɹ�d;~d���j�e�a��Ld`y8w�/��W/��Bl(h����ū�&�ATA(}�W܈��MIpT�>���m�uq� �l�^����R(]|��ݮ���i��Z��x�j6�j�L*�~��
�d�ꀯ�H��nq�G_2=_�螄�� ѕ7x.C��nyq$�R� �Uv�=eHF��cE�9)Q���m�M��&^^G���"�W#-5��x}=c��5X:7v$ԥ�>�,~Q4-#n�i۞�l��+X:TV<�ѣ8�xI��ε� ��Hr�3F�S��5���B������uQU6��Q����9"H�Zzk���l] ����4�K*n$��fg]:�%��ɹ�]X�Y�e�l^7}������hU�f�{�=�
M�r��^k,�^��5yn징k�Y������^���9�v�x7�~T�g����ʫ��n���p_�ʐyZ�� =��P{uz�6L�)�E8�����+� �^�h������j�UOs�R��t	�Y�\�J
����a� Gˊy��Q�xqq`I�~ 4&´���#�k>�M#6�Wb"w�����ڟ�VP�f+��h�1ֆ��������'Wy�6P�ei��Y0���w��L��@��ѱ0O��(z�p@U���`
��G~�Ӧ����pI�R
�f��F-��T�<�a:2%�^����4��
j�BP<�����=�&�W�������tn���y���1Ƌ�QF��_��.�8�s*_�՛�r��w�JG��Պ|g���+9ho�����9�ۙ��V@�fz��ȯ��u�}����Xq/k-���:q6M�H�欨�0R�T��q	�M�xf"���t��
.�B������/�*Q3����cẋ�dN���K�ǽS�bkFT^���"˼�����!kY]sQ�O����?s�r�U�G�a��2�^��ߥٹ���D�����f�p�ƌ7z^��$s$U���s�sfW�Y�+�X٫����?�SxN�;�� �%�L���yrny�e����`YNZ"�Ҁ�>�TEp��,��f�1N���DR�sD_~b�]�Q�|�`�6�+��bF���+kk���o�FV.��%9��7��}�G��n9q��@4.�}i�ܾ����z+l6E}��`_�,���V�q�o�up�e�� `�U<A��!?�P��tUe��u3?�q�"ʭJ®���@�TP2�s-p���,�O�VV�}�k�d��I;r�u���eOCơ���]�1��3rZ�l����q^$��Ǖ�r��D9�׭<EH��c�����'Mm�5^w��2�����}P#=l�1��I}�����꧵S����-M�d��͡�2�� øL:!�H!P���@ټ��ru}���:��S�s?��t�X��둧�bC=D|�5U��~��b����IH/��Ϋ>ݷ����Kc �J� �<�j⾔"�f~̑Iuҗ����C���"թL�C�_�LZ@�����זxf���(�В.�y;g&Д����P�2��H;�N��wQ].���t����J��XE܇���SRT�Z�j���ˮ�M!o!� cLS
U"~u�P�N�˻q��%o�~�"�a�����[�:�o��=�i=u��2�lHH'*�����͙��ï�w��H�3��c'Q7݉��������m��6���K��G{aK�(d��R�w�=��?�_�G���X��� ��Ǐ�&�' �5)����ߠ�œ�	�Q1u-\�5���x������������F���/hʤö��~ʉY��k��D�~� ��,F#N���Eĵ�����|X�=ԁ��'%ѝA�A��m�Ч��[�l^� ⷱ�����/��/K[��_I(��/���U)�Q���2w�y��mr�z�Jc��i�W�o����o��Z��fO�oi�6* ̳3Z�|��Ɩ��I�/���������4gt�S���~�aɒxn�6A����V��5S�5�=ZeC�1�W�S��ly�(���Z��K�r�N�C��2$��"}�g�F���N�u�hI��UZT�Ǘ���QJdgl�3���Z�l̐���&��U��?x��|���@��L+�U[�	P�i�U���Y�ݧKG��̡c��K���"��
�q�m'�T+���}����{��TY�3���/�z�Ș�>�E�"i.�z��w�����cW�1�o���ݴ�r�9�6�.?8���Me��*���?{A�E��c�bL
n��y��w�Jp���Խ�O��̷���X�����������#�T�5FP��b�����N�gO=3��+.�5��;�>��rɿ����=���'����H@��}N��U��3vտ�,�M�oTK�cX��VU�i����X�?0z@U!S+X���Зm���i k���O�Əzy6�x�",�XJWuU(�/S�����fM��F�������܌6�m�/(�n�Ѽ�ĉׂ�	�1��cf4D�#�6�lͫ���L���l�|E�
\R|�=珿_�Æ?1X�V(V�%7n�zح�*F�6@-�'�o��������*�����R�bϸ�j�Y/!ojݵgl�[�*E�
 ��Х0/��A���'Kd�+���^�,�_��0v����w�_�˝���~!�`�u~餍�s��x[�v{�Y�۟�8� �z�����MY�k��#Z�Wr�������N�vS�4���drI������Wh�,��ԋ�X�E�U3�8@������%2+�j���%������n��[)���+�Kǁ��3q �?��^֟u��N�S�N�Y�Ð�\�"��RQ׋�['��#�1��^�r���(�z�I�]i���4;2��ʙB��1p��[�Qno
 Q�+��u7Q|}g��lG� l�=������Ce?��޳@"_�L��X�l~~���Y5����?h�D���bD���U�a	��3��-��ۥld�gH��r�ޤč}�F���.�Q��E�i+$?��'r>��i�}�_׹b��Y�V�v�s����_�nk�J"#�N{h�{7}u!�����n��R3�s=|����/��s�˩@^7M����=��=x�級̢��a�{�.R'ٝ[ً!�!�L1�(�z��$z�����]����*�&��ŉ�T���1��N�3n���c����$�@��;�-��=�q�x�#�:^1�� �T�_�%`o}��?�����&2�}��:�5=����:4?�&���Z�&����:S�,2-d ��퓼Ɋ��р�JU���[!���{�'�gM��2��Z�}Kr���9��]�P�9��Ac���P�S��#�u�n^��sN*���à^���7�	ߕ�p>�l}�ӂ���Z'R�y��E�e�/'b�%@��3��Z���
��.����V�A�H�K-O����Õ�n]�it����6 ʆ�7Bo�'� �5H�vl�K�F��=Ԍn �F�c�i���̎~\���3�/"Z-���8��3p�z�}(�L�"|tYz~����?Kj`g�ע�		�
�x{��;s�$u9�+�Ĝ��|���}�]�
���׵X14�9�KO�E��=��?w���p�9�{i�ks���oip���Ww\�\��{�"XA=-c�b>����ǈi�����f�ǜ0:���sh�;����QC|+�U ���B��	��O���H\a'�N9%�[��c`n�c�N�rn�����۞��:�f�h�n�[vZ�_�)r�ۚ/1����S�í*	���W���hp͕�?�z­�����8ڸlx��d�i�:��/���zE���PK   .{�X6e�b�  �  /   images/c0cd0a79-4e96-4647-8bb3-400a2b193618.png�YePЦ=�8����<Z���n$D���H�n��n��n	ii%�������ogvwf��g��_;��j
�x4xhhh��Y���wp�Ÿx|�	�a����������h�+R���k;Y�{��Z�yyy��stp�0s�z��j�y"A��F�(+����7�R���4�����j�����0���Ā���K���%h+˻���#�����SH�L"��8:c��X�d��˦��~����F'O�絍׌��~W��z�7|��;����d�CD(�Gg����Ȅ����S`s[ �OME��%��!�HK�VP�'�M����<���fU�*6��(�1��LH����u>'��?A��3, K/56���'���W�er`	�<5�WåvR���,�Du�b%�\Β�Q"G�Ni�p~ⷄ/��0Z�a���3Q%�`>x9�e�1#�b-�X��,�Mp� /�ɝ��� K�C/�*����&�U���oґ�9�N�#\������;ɼw֠u�PO.�s�V�q�K��= O�}�)(IH(q77��En�3���&���Z����[��n�:�9��İ������XYܞإ.#S��(CR2��Z�V�BXp�Ll�#M]���a�
�-f�*�&�үN+6h2l��Vb��9�"�%��Iʿ8�}NFA��友_p�V$�n�-B=���į+�����"��>aH5ğ����i����V�:ܞMpi�/�%�������0�Bh�I�e�uv�8��y��.*M����p��v�Bf@ 4�۶��u�uR0�f�JQ� ��Ǵ����\fZ^�9���7���#ps�:�֮F��*�+���g�M��}��D,H�����Y������W��;����y���#4j�}����>���˶�Z��g�K��h���Rǝ�}��dp~	�Z���=�)f�9��F-�g>iCb�4&!������&�ֽ2�����v�
��&)��l���&�(�	����ƯVjzo��2���{�����)Q�z����e�GU�����nS�US����6y�j�h������#k�EY�AE:r#��N������&h�U���q-�^⑼���ԛ����ԅ��I����~(���Q�T� e��0��Y�5�V�1�B�F�mo..ݍ����#;���>*��Td�rb�}鯻|��~J�擕�,��\U�P"^N������wT߶
�����R@�����9�b��u�pޓj+�|}�=����W/d��n��2os.�E
�k=+Z��#dK��)��m�L��<�a��gI���*^�"��R<��':�`���U����/B���տxNsW���U�N>�x˒�7��I8T�\#��5Q��p�g�4�~β|}������+�n� L��΅�?^CV��r�q*���6�Ⱥ_r��4��ѫ]�jIV�9������B}�((�������w;Z�ƋJF8��M�S[�Z�b��������,����Ju��=�a��,���ŬD���^-[�9�[�u��]�ҏ⫃�"���G��er1��&e��.,xí9�z
q��h�ɰ�i<�G ��0����t�/w"m?`M�,�m+����T*J�]N��_��fw�^{u��|o>vO#���j��Lg8���d2�&�Z��b�؍0V���f4 �~�h/ͤ��
_�{� ��A�I�9y�����B�K��L���<b��o����^ZEC���`�a���?X�5צ����b��K>�3&�.�
k��C�K�=��Pּ̑��j��a�RqF.�ZFЖ�-�ΦnZ��v��*zy�ag/b���@z(����l(����L�R�E�8�7Ȗ��f�0�9�nk\����5=^�����>uG_���?y<nP�@5�9����jw��>���a�6�Z$�?2�ß0��u�qB����;��x�$�8��.�sFy#��Z�C�z��R�
��m�#B�C���/�p�!� �p��c��kbdl^Ϭ�'�h�u����@w��G��q,�r���5��6,5R�w��������!A���Irܯc��A�_��y��n���1+�2��"�C��Pb݀#m���`�|�Hf�����F M�c�7vQ���ݏ�I/"C��Qc�3v:�J��:���j����B G?L{�hP�S�9,�oc
����w�B��/3�������J�ˉ���l&W\`�={�'
���]Mc���H�Z���p�OI�F�ۇ�[2�)��u
���&D��x#l����Gq�!*)/�*�qK�I��*lq��^��{数s*G�MRϿ�?4���(���@rs�s��]l���f�Xy��c�R�F�������SiC�f#�?2ښiZ [�,�9+�$jw��i������LV�	ܜ��'E�
�v�!"��o��}*<�Z>Z���0�l���2#	O�E�}H��d��
ta}�����	�����p��j8�����έ�8�4��'"��Ӷ#'�zT�!xY�6N�,n�1^PL��]���}��\�����1��)����m[�T��N[3 f'�2��[��:��S!���`%ۢ����"���"b؄�����"��=�N�BC��@�%A5C�:�����n�Z{�qM���?�2�Q/:j,|�w�f�6�.�-�f����l���:Sh���E���K�fg%�A��y�^ǔN�e�������U�k~��0�9�1�x�\pѤ�y/�Q�\2M�yrn��X�!�xG$=��hm/�`^V���Оq�w}��#Ǘ�M
Q�.���u�+]>��GQW"����SӐ/�!)b�|�n�ʹ���^�T�D�@��s�D;�sN��L ��s������hHA����r�N�u"VN ��9$����O�����x=l�f�X�I�8fWē�[�|�����Q��V�bl��%�`��������Y�&��4aon�*�՟|F�Q}�~L�o+���_R�#��'Ҹ&��-�#���L���'�����fW��ķ�!G�4bK�8Y-D~z]�v ����Y�ˆ�;�=^�װ�����<��n{�)n����BI�)���ltm�{���&'&|kӛ|�~1��3g<�
Aʈ%afs����$$xHl7��|:R������FY�6Qu��)���ӡ죢l>:��*4��?�bXcF�86ԏq_Q��J�KZݍs_Yg�_\��N�.����\�;�����-)���Wn��M��lgӠDjVT.�痏RěA��mk=�������T��>��oE�U'�6�ȖCLn�Jy�辶� ���� 	ө��a�[�[��?.�=�s�mp#��~�n��io���٣���m8�9Ɇ�GMD���79
&�ۢ���,0!Gl�ݝ^3ɕ'h�����]�����'x�
,�Uܕ7ě�w�wr�!�ڌ����z{q�\^X��Y�E��ދ;��[�p!m�����}�9��ˈ�6D�7��E��_����A��.M�p~�ap�~$�S̲���2W�}�7�X<6v5k��w6g�&����/��H��leIHzj)�Lt�fr�ۙ�ͭ#�+�o��������kԏ_����k��S���I�� �lVл~�>��Ͼ�]��疽�/��m�x��7=������>�-�dB8F��*�]� G������șUIT�1c��'>���������f4�fq9	��s�ҿ��d݂�)���]y�ELf:���(���tP�����gn8�}}S_u�JϘr��|�=\�P���r�oRE�Mo�pmm��<f��L��'�g;� _QSc�v���TFbX��G���ݾ���3[��w
���V�����j}"5�d��`9�x�&���Ϫ҂�j�i�S��_S� �g��b#.����!����Dy�9�rnyԶOZ�����;K,gR�2�T7�,���o���RHQd;���%��l`��z���vZ�ɴ�J>��#J�*�v)s5�[��o7P��
uޮƺ�f�pk	��{��;�Q�TR���(@������ę�w<���њO�o0-ȁp��÷���$��Φ��0�J(���ګ��z��/9�nD�_�j`:� �b�j��3h>y�5E�D��2Me7�.��np��ޱK���I�u��{[5)����J��}��O��-b������&C�I	���%�)��jן�\o4�1<Rj= ������z����K�L���uH믒�"�^�g� S.�T� 1|V����!LPv�!��$[ 	�������Tsy��WKvJ<�aXv#�I�t�H���`F�[Qz��E�n��`�L���m��PN�AAQ>�"���`Ѳ���36��ˏ>���f��d}j@�D'{�/h<�c}��s>�q�/�6�Q�:_�����df_���������P�&�:4��g#�����zx�(�>ҥ�X�w|����|(�"���*���R�g̛�>J�B�Ok�oD!�mH,�/fW:X�^g/!���]w��-wT���Jn�}Ja��2�~�f<����:����,�F�w����c�-�Ѩ;���*���s�ڴWf�zC�!�oQ~9��(����Wc�>�9Ue��T�%l
���M� +�R/��f���#��|oÈ����@��w:%FEi9�=�u���c�ceh�����g�9�������F5�p ��5ony��Ċ�ƑX� �I?��Y��<�M��O����˺OO|���N�9a�-�q�0��Q�ͦ�+[�k���1�����i������=۪m��M{)͵�uV�7Ƌd
�*8�hF%p�!�Y����V���Y9�)�����7���]��ޛ�ݮ0�"�0�΅p�z�R��l��+�Y�>����3W�D�����Q#�Z��e��i�05�Ԛ�ì9�� �R��������{1iR�8�wy�'�'��8�
�DX���A4_M�;�S�h��QY��}�e�#��-�m�X�!�V۶
��1�M���*Hj;�D������KB�O��S8i?%߼��MRZ��m�E�q�`ʣ\m�K�#>?v�[�Ռg-E�{f|%w9�8Fu�ű�����K�� ���c�����J�xhM]�e�:F��G�1HL>o���c6���e���a�{��aKL���鹲�Ap��8eo�� �������]-���Td 8o�{��M���q�c������-�p Xp�Lp���~&��ʭ�Q:psk�����c�Ui�/c��$KQ`�x�B���ϟ��?�:�8���܍��>����<��� ��$�Ga��D��O+������WSD�,��lCNP���6�7�ȏv���L��P����gxE&%���������S0zS�)k�%em3�
���M3�z��[�ī3�r���{l��1���hp��ՙ��d:���j7����9-�C�"�Χd���eߣ�z�If&0�\�/>c�BW��|P�x�Y�[(ɕ��H^�?���	�M'�������7?%ݽ�j�3-iW7}wX�z�.KP��{@�t�[�QC��I����,d�<r��i�7^Hkɹ�>0ا��ȫs_&*�~�ZQ���־�����=>�z����*w "r/`�=_��?�}��l]�R{i�x;Q����4J�Z���3\�����jh(!����K���x��
I������\޼� 0��+���	t�$�#?BzF`��3p݀��o2TT���$pKt�&�a�
g]�-W$.�����Yv��G�����������0������|d�qS�E4╬�3⓱6�ڒ�=���:j0~�l�O-m�C����ҺQ��*VZ��n�'�FQ{���\ld�B�ȱ��Q�:��+KT~�*����?�w��lN�:�c�Dh��Y����y�J����,$���Ǔ}`�~�������C;찤Ƕ�#�l#��&
�{����k���%��N"���}cf�df.�,�K��#�>�g`Fv4�O��9��x�9����?�6�?0o=;R��L@�����������?=�Q�a�k���fF����3GТ�r_�������@��:�u'��"��+?ʳb��x�'������#����C�a����e������}p����$���͍��&N���v���s�;H����$(��贒!�������FŬ����`V	l�K�5V��� 4X�G.~'�:��H,�9�&{�5��L$U��m���3M���빮�;��I��y���I���[}��1���;@���#Z�
���b�@�8��J{��=.�Ѣb�.G�+���_HiIܸ9�fqe�O�ߣr'qx�0)�p5�ʒD���¹�Ⰹë�Oqp��c�U3��Re�F..���ߐ��k��/�0	V�Jּ�l��~i<\��̼E�paTT`�L���W�
 ߞ��YK�_K�Ǣq�S���SI��a�\�,t"������e�ƪ�jGTNG`����˫�7B�Γgh��\'F&�^�/�D��˽��%5+�GE�B5tM�'���a�GXh'��s����՚(pFZ�I����e��0m�������?7���M�⛿���;#cU���[E�z���D9#t�1>��;�o[]�=�Rн�G��02�3P�`Dh�v��f=�Nl�:�^g2�������:�:������S`���g*w>I�%_����3`��RO���*�cl~���ơ��}إ��閍N�eg{J��N��Q_3~3�[��`���8���@i�";��h�q�Oov�:�_i���m͉C�k%�w��ǹ�&J���]W��k��b|��#� ���ny�� H��];.�
	��;|�}�eڽ��vV$�&������H��UĮ��c��8ꡌ�ߥ��GZ|� �*ז�N�)*�j�"'�DI��!t��/��Ƽl1�#��j�(��ي�ǧ��iY0]|I��C�#���}������;?b�(���r��̊��~(M����G����W�Ȉ��N�2�?��e:u���9H���E�u�ƲGO�_�1NV]��^$P	�7�[y J�Fb�(Z��Gh���� �d�W���-��A�Z�Їe��G�>��Vϰ����C��h�^��1q�%փq�5񣅨�����a A�9�jl��tflR���b����+9I�3� 	�$_�b�2ػ����M��Ӊ����wK�i<��7�~��yɜKR�G�1| 6�P��ҪotF��TPS��P�ӌ��C	!��i����D�X��y��>��M��ߋ�h�U"�,z���򭁏&�=U������.�2���AW�Ԗ�g�՘����<5w��i�\��H���6����?�?S�S������PK   .{�X/yR�c  ^  /   images/d2af519c-c065-45b5-bffd-6bf239de2b90.png^��PNG

   IHDR   d   P   �	��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l��gw��c};��ΈU��ф#H�4�� �U�R����HU�V�z� �rD4��F��\���І�p8�Rb0�41���X������lf{vv����>�g��f�����������*�8ˏY&�d�xY���/�m\�BQ�6��#���a< )���������������~��f���rݟ���M�s���Ȳ���x= �IaB�� Zl�ۗ��������p�I���zV��ˊ������۷��v��/����,���$1�#L[ 	����t�ҥK���_����Y@NN�;wn�RRR�_s�â�Ͳ�e�[,>�7�AI�5DĐ�ˢ����I�&��2�M��	b���j����͇��cg��3,����r�x@c�0!W�\�[vG�p8���/���#�)��Qr��>��3L�9�e�OX6�FN�^(�1G����:joooHKK���"����.ܻ�e1�wYv��(�S/��t����P�������;D\I�Y��;,+YvRT���h�p�Ȼ�������Ғ3x�`b����M	��*�?�4�@�!�R�?x;��������/4A>��E�Yǲ�4W�{��(�ۉ	2n�8:~��~XŁ�Q��UWW�C��������Y^e��
&c�MFyy9�]��� e޼yqՏ�#)S��kg%���㏗s�=m���Ɋ+����
?o.?g3s��qLA��À�"V�k_�n]\�8�OI	���a��ڵk�9+2d9�N�&�|ʔ)t���)��@��<�zۇd)R�)���d�x���F�O��dgg��W2�T[[K���b�-�b�O�>B`�[�{������p�}RC&�6�gXo{�!��
b6o�L'N�S�N�p�]�}���Ni1w-�u ��ѣ�\�������h�ر4|�p��ʢ�S�Ү]���=�R��`8�)1���㡊�
�Ng�QSSC^�W([|���)4!H�"�T��u��bK�)wYY� %�� ���w������1		qdCo�B�p��R���L�'O�dXq;x�~��i6l�p�S���t����DEU#�)���y�2��SK��י �`\o���bU��1���@q� �Sc�����̌���A�Pt�K���7n�nJ�S ��Յb��[dS��o��f�q�V�Q��2(���]l}�4Q_?F�~l��=�������F���u8�)ܛ����R�2-�W�^d���is�uD�NXCC��5e6�u�LG+=9t�;؅����j������)/�y}����D�?蠃��G��M�L{��P�/�f�Iv[����-���p��N+�n A�&��y+')A�ج]J_�p�-�c\	N
̘1��/_N�������e��	VBA.�qd�̙��~I)h�v% [�Jo_�25ys�R���ug;=��h�����=[(1\���TO-���������tQ/+��2���Y�q,��!���l�U�������dy��V�WLt9����'��IA�0`�Ha�]�d	m߾�������`�cdn/��M�0!|��W�
f$�G�|���B�����a�r��.QN���E��S�e�l�t�(��9?�f�n$���,��4�jNO��"t$-�����A
Z<�pa�c�ܹsE9b\Z=������D2n��Ѱ���RЪ�����\A{/L�*�B߻<>l!�*զ)��qd�����.�a�7wO��n�f�=�<����nR'F���@�$��R��"�����/:yP<�-V�.�0ta �3���j-]����nѢ�lXHt�bq�C5����
�B�c�X݋Z|Y�V�T�����3�x� @]){��$�]`�� ��E"CF�v���`�޹�yp[pu�`�)�6�:�.�f����.�d@y(3[Ay�禋Q'��]U_	i�aAqA��ߣ�=�v~83"�{�V�,��1	]�p9P0������"�Bl!dVp] ���*�!��9���6_F�֔��Q�^�}(<�Z(�X'\n8}M��(
�Ҭ�4��2a!p;��mA�1z��gg �
��X#�fʰZ�Y�xϛ���1	ٸq#Z��髊1&��D�(n1&V�n��L�����Q���ƾUg�I��Ç�Q0��p�BJ��;!2�����X �C�Dn��ʕ+A�ZZZ�$J���28�T�y�f�}�>~ժUaRt%n0��TX�c<^!�,�IQ�u�����%�@�#�MT� ˈ�E'����6�=��z��B0�٤�H�L�w����!��	h����A���'�ǃ�	��SIH$�	뉢����!	��A�9�SS̰x�bw�@�u�������8����.��$���Y�9s����e˖)2�Jʃ>�zNN�M��֬"yܬHH�oD�F(�E�`�A[˒��e@�1;(1	n�[E�#�$����4���0xXPP�̟?_]�z���z%)2�?�p�\J�\��G��`���eI��X ����;��Z�;�x!ř� eŊ����ۡ[�СC�"p��c�xԨQʢE��M�6��d�HpV*^�q�UB?7�|������*���4�u$?PLՑ����<v��1hXb�q�̙1�����o�6��i)=�f�4к�:����yx?oڂ�0�����{����z<�=�-2#\�F�H�{���z	�~l����gY���O��h�uf0c�����>eVl}>�d��K�,ccU��P?z��k�Neǉ'�<�	E2vt����Ԏ��[�n5�V��$!�!:
����$B�/	I!��=ѧJY�"m9^,�!	Ijk{y��?��Kښa/��.*bJ�$$EX�tӫ���XxlK�dXb����t30��fڲs�ӣ�ZX�f	o�MZ/^ZH�C���늟���w�ÂD��&��$����38�MXXC��XK{5bU��O�諟It'0�T�vMu0Ȫ X����/�~¿"��t;LQ��'+}ݠ|>5�4��e?�v�߰%���?|饗���nX��,"-��;8��,{YvKBR��_+��wi.��1b�|IH
�ي��������_=�3�A��,��|��Q�\IH7C�)��+W�~��XO�e&��4ik�1�=����nF�UX�h�ol#�k��W�he�g����-$`��0���RFZF��F�e-���PW�`�ΨQ�^����>Â5��(�|6*<,	I�m�ǌ�>��e�|������,��V����ǉ�H�B���z�����_��V�B�0�.�|�4��$|��9IH
�q!n|���k�}bj�UB���9�X��]g�0�����V	��=�Y��D"��Κ�7�,dYb�|����$)�d@wm�����0)O��)B��fA���u�u��l��"��`���N���x�]?�~���&�e�_w:�x�$$�|��#G�|�ԩSq������A8c    IEND�B`�PK   .{�X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   �|�XLB�}�	  S     jsons/user_defined.json�\�n�F~A@��a�~�?�Jw�u.��l��Q����&UJJy�}�}�J�/�H�Yw-�(�s��|��8�e�����z�_|��<��d�1��y��(CN�,׶j����������}u�a��j��*\���j�s��n /&�Omc��8)@���Y�A3@c��<(B*��zQ�!_��9�'wxG�rn����+����;o��]:�I����=)��G����L��]�o/��+���m��::

�kA8��J����\��"ž��>^������<��b|�e���g����|>)�RO���eB�fw�ΊO�s8�D1�����:���NQ�/��������ye���*}C�ΘbBO4�K�����4w�2]��+cCu�_^��_'��q��G᣹Z��wr҈OZܗ����Fx��~g��W����}ѱ{�O�ֈ�[�������F�% �����׍dK]�8K�"���էy�T�k��,�\�7�tQ9�P�N�ώFo?��;�>]�øY66���{N���I�1���w�`�'u�׫�zU������iM��`
��$F�0>(��#�N�l�_>T�G`�2��̓nN��$Bh�$���Z��7��p���Y�T��?>���_p2T��:sרٛ��0�ƙ�I][I���萴�q���~B]��
�������m�	n�X׋�*��j]�����RTr��euS�>�^�'���z^%Ȼ�r^��}W��֛|�tvյM6M��ƭ�e(�?.�S�|��k�1�"#`$�J�BiPX{�S�x��v[a|��6��8U�P�`�2F��(	*"*��.��v��Zw�C$�#��Xkc�ڔ�U��T�K<���k��9J�D�`)l�@c�����6�a��䗏S�c�D$��!XU�㸤>�(���2U�(��1� ӣ{�ʦv��@�?*egl3��Ӑ5�##u⩮�+Ku�Z�
2�bMV�Y/��G��Ƹ��@�qn�R�)�9�#��v�zA�Ou\`��i�6�v��Gè��\�cr���ݟ���ND0 �4��t�iS�Tf�&�h�}:����|�*�=n�erf7�&I�r�
�1�9�^XS��N9nZ��IWPÜF �MRd+(�	�ZD��	���Kz&7\��R ���04��{ӳ�+�{����
9L΃����uu����1�w� ��'���=Vl��!6W��Y�T���I����'}r���;�o��P>�;�ߥ�b�y��c���W(���6G�Ϥ�g{���� s��ͫ����u��/�|��b>�l=T�t�> 
<}�2̂��c$	��	����"�0( �"�0( �"�0(B�"���c�k�n�Lb�@m$���@M@�@R!�"R]5����(NB��D`)���i�O3ɇ1������"��MSk��,��`y׬E.s�[0�ƕ+X���}�M��I�G�Z_�9�1:��};������b�+��R*�a�k��;�xb"�ځC�㖃�уH�I���h�=�0Uy��R������T�����Ο��Š�Zj1�Š�Zj1�Š�Zj1�Š�Zj1�Š�Zj1�Š�i����2��h����HweUWW)�6�@��tc"��4*	p]�]-ҝ�C���G�Q
�E4&
$	$jM��Q�o�B0� ����(�rOWjY*�g�Iƽ��t9�����_Sg����=����=n�г�f����[|������=V���n�mK��k�o�I��!=߂��Ǣ�[p���XP���y#�j�V�E#�nĖ�e3������}p��LӮ,�����H�Y
����	:��Y�z�LӮ,��Y�z\'�xT���`xѼ���U���=$�O+ĸN\�W���f�:wE_-�6����+���YxH����O�5��,z*�Y�I����&O���W�T�is�%-��H�i�h���I;mVN��َ���=�����	Kߵ���v�e��mkZg-���Ī���$���>���7͆��sW�Nb��d������e��~�7��
�����}��-Y������*�mv�?��´r�_�n��O3�p7C��Վ!��u�p��� )��1L�O�^&&�F�f�
������|���Lě�Ӂ����z��R��AFAnvf��qJH�1��}��Ѽ5�
.
�Z
&D�#❰�����U�<C�Ѓ{��Q���?݀%����	V�f�JEۧ��t�ؠs�Z����c����g���`I=0n���L��,���F,��p�^rr��]�O�|ħ����x�~���n�r~<��Osq�C�<����H��f�*�0!`�b�<C*0#�/��4zP�D@�+�Ml'��L*���2)�=�g�1�i���(�2��f`ڒf۟F?�ȶ{FDeD�G���JsN�3�2�:��9������H�E��F�@�6�?y���xA�o��q�Z�#������|��?PK
   �|�X_�ά9=  m8                  cirkitFile.jsonPK
   .{�Xh��;�� �0 /             f=  images/08e4a639-d7b6-43fd-85af-03d86c8bfac2.pngPK
   .{�Xo�>��q  �q  /             ^, images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK
   .{�Xv��� f~ /             u� images/4d249bba-3190-4770-b321-fb8fc027a237.pngPK
   u�XY�\HJ  �  /             ��	 images/57470e45-49b8-4c21-99d3-774ad112c262.jpgPK
   D�X�Rr5�  5 /             �	 images/5dbae223-cfe3-43b3-aef6-7502dc6b2367.pngPK
   D�X�@M��  2�  /             �Y
 images/5f70de14-173d-45a7-8b46-cd4e4e8c904e.pngPK
   .{�X��p� �� /             ��
 images/7e81f6ad-0912-4ff6-bfc6-e58bb7840941.pngPK
   .{�Xd��  �   /             �� images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   .{�X�r�44  /4  /             � images/863c2d63-52da-45ba-83bb-7a6a6689309e.pngPK
   .{�X�1.:�  )  /             � images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   .{�XN�v4	� m� /             �! images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK
   .{�X?S��� 2� /             � images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   .{�X	��#u } /             � images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   .{�X$�8�l  �  /             Y' images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   .{�X+L$��� �� /             E images/aad47697-5cf4-402f-a095-abba84463b41.pngPK
   u�X]��  A  /             4 images/bad899ba-ddb5-43c6-9f63-2d962537fb78.jpgPK
   .{�X����<  �  /             n5 images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.pngPK
   .{�X6e�b�  �  /             �S images/c0cd0a79-4e96-4647-8bb3-400a2b193618.pngPK
   .{�X/yR�c  ^  /             �q images/d2af519c-c065-45b5-bffd-6bf239de2b90.pngPK
   .{�X�GDU7� �� /             �� images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   �|�XLB�}�	  S               	d jsons/user_defined.jsonPK      �  #n   